* SPICE3 file created from sky130_inv.ext - technology: sky130A

.option scale=10m

M1000 Y A VGND VGND nshort w=35 l=23
+  ad=1.435n pd=0.152m as=1.365n ps=0.148m
M1001 Y A VPWR VPWR pshort w=37 l=23
+  ad=1.443n pd=0.152m as=1.517n ps=0.156m
C0 VPWR A 0.077431f
C1 VPWR Y 0.11654f
C2 Y A 0.075353f
C3 Y VGND 0.279009f
C4 A VGND 0.45021f
C5 VPWR VGND 0.781009f
