module picorv32a (clk,
    mem_instr,
    mem_la_read,
    mem_la_write,
    mem_ready,
    mem_valid,
    pcpi_ready,
    pcpi_valid,
    pcpi_wait,
    pcpi_wr,
    resetn,
    trace_valid,
    trap,
    eoi,
    irq,
    mem_addr,
    mem_la_addr,
    mem_la_wdata,
    mem_la_wstrb,
    mem_rdata,
    mem_wdata,
    mem_wstrb,
    pcpi_insn,
    pcpi_rd,
    pcpi_rs1,
    pcpi_rs2,
    trace_data);
 input clk;
 output mem_instr;
 output mem_la_read;
 output mem_la_write;
 input mem_ready;
 output mem_valid;
 input pcpi_ready;
 output pcpi_valid;
 input pcpi_wait;
 input pcpi_wr;
 input resetn;
 output trace_valid;
 output trap;
 output [31:0] eoi;
 input [31:0] irq;
 output [31:0] mem_addr;
 output [31:0] mem_la_addr;
 output [31:0] mem_la_wdata;
 output [3:0] mem_la_wstrb;
 input [31:0] mem_rdata;
 output [31:0] mem_wdata;
 output [3:0] mem_wstrb;
 output [31:0] pcpi_insn;
 input [31:0] pcpi_rd;
 output [31:0] pcpi_rs1;
 output [31:0] pcpi_rs2;
 output [35:0] trace_data;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire \alu_add_sub[0] ;
 wire \alu_add_sub[10] ;
 wire \alu_add_sub[11] ;
 wire \alu_add_sub[12] ;
 wire \alu_add_sub[13] ;
 wire \alu_add_sub[14] ;
 wire \alu_add_sub[15] ;
 wire \alu_add_sub[16] ;
 wire \alu_add_sub[17] ;
 wire \alu_add_sub[18] ;
 wire \alu_add_sub[19] ;
 wire \alu_add_sub[1] ;
 wire \alu_add_sub[20] ;
 wire \alu_add_sub[21] ;
 wire \alu_add_sub[22] ;
 wire \alu_add_sub[23] ;
 wire \alu_add_sub[24] ;
 wire \alu_add_sub[25] ;
 wire \alu_add_sub[26] ;
 wire \alu_add_sub[27] ;
 wire \alu_add_sub[28] ;
 wire \alu_add_sub[29] ;
 wire \alu_add_sub[2] ;
 wire \alu_add_sub[30] ;
 wire \alu_add_sub[31] ;
 wire \alu_add_sub[3] ;
 wire \alu_add_sub[4] ;
 wire \alu_add_sub[5] ;
 wire \alu_add_sub[6] ;
 wire \alu_add_sub[7] ;
 wire \alu_add_sub[8] ;
 wire \alu_add_sub[9] ;
 wire alu_eq;
 wire alu_lts;
 wire alu_ltu;
 wire \alu_out[0] ;
 wire \alu_out[10] ;
 wire \alu_out[11] ;
 wire \alu_out[12] ;
 wire \alu_out[13] ;
 wire \alu_out[14] ;
 wire \alu_out[15] ;
 wire \alu_out[16] ;
 wire \alu_out[17] ;
 wire \alu_out[18] ;
 wire \alu_out[19] ;
 wire \alu_out[1] ;
 wire \alu_out[20] ;
 wire \alu_out[21] ;
 wire \alu_out[22] ;
 wire \alu_out[23] ;
 wire \alu_out[24] ;
 wire \alu_out[25] ;
 wire \alu_out[26] ;
 wire \alu_out[27] ;
 wire \alu_out[28] ;
 wire \alu_out[29] ;
 wire \alu_out[2] ;
 wire \alu_out[30] ;
 wire \alu_out[31] ;
 wire \alu_out[3] ;
 wire \alu_out[4] ;
 wire \alu_out[5] ;
 wire \alu_out[6] ;
 wire \alu_out[7] ;
 wire \alu_out[8] ;
 wire \alu_out[9] ;
 wire \alu_out_q[0] ;
 wire \alu_out_q[10] ;
 wire \alu_out_q[11] ;
 wire \alu_out_q[12] ;
 wire \alu_out_q[13] ;
 wire \alu_out_q[14] ;
 wire \alu_out_q[15] ;
 wire \alu_out_q[16] ;
 wire \alu_out_q[17] ;
 wire \alu_out_q[18] ;
 wire \alu_out_q[19] ;
 wire \alu_out_q[1] ;
 wire \alu_out_q[20] ;
 wire \alu_out_q[21] ;
 wire \alu_out_q[22] ;
 wire \alu_out_q[23] ;
 wire \alu_out_q[24] ;
 wire \alu_out_q[25] ;
 wire \alu_out_q[26] ;
 wire \alu_out_q[27] ;
 wire \alu_out_q[28] ;
 wire \alu_out_q[29] ;
 wire \alu_out_q[2] ;
 wire \alu_out_q[30] ;
 wire \alu_out_q[31] ;
 wire \alu_out_q[3] ;
 wire \alu_out_q[4] ;
 wire \alu_out_q[5] ;
 wire \alu_out_q[6] ;
 wire \alu_out_q[7] ;
 wire \alu_out_q[8] ;
 wire \alu_out_q[9] ;
 wire \alu_shl[0] ;
 wire \alu_shl[10] ;
 wire \alu_shl[11] ;
 wire \alu_shl[12] ;
 wire \alu_shl[13] ;
 wire \alu_shl[14] ;
 wire \alu_shl[15] ;
 wire \alu_shl[16] ;
 wire \alu_shl[17] ;
 wire \alu_shl[18] ;
 wire \alu_shl[19] ;
 wire \alu_shl[1] ;
 wire \alu_shl[20] ;
 wire \alu_shl[21] ;
 wire \alu_shl[22] ;
 wire \alu_shl[23] ;
 wire \alu_shl[24] ;
 wire \alu_shl[25] ;
 wire \alu_shl[26] ;
 wire \alu_shl[27] ;
 wire \alu_shl[28] ;
 wire \alu_shl[29] ;
 wire \alu_shl[2] ;
 wire \alu_shl[30] ;
 wire \alu_shl[31] ;
 wire \alu_shl[3] ;
 wire \alu_shl[4] ;
 wire \alu_shl[5] ;
 wire \alu_shl[6] ;
 wire \alu_shl[7] ;
 wire \alu_shl[8] ;
 wire \alu_shl[9] ;
 wire \alu_shr[0] ;
 wire \alu_shr[10] ;
 wire \alu_shr[11] ;
 wire \alu_shr[12] ;
 wire \alu_shr[13] ;
 wire \alu_shr[14] ;
 wire \alu_shr[15] ;
 wire \alu_shr[16] ;
 wire \alu_shr[17] ;
 wire \alu_shr[18] ;
 wire \alu_shr[19] ;
 wire \alu_shr[1] ;
 wire \alu_shr[20] ;
 wire \alu_shr[21] ;
 wire \alu_shr[22] ;
 wire \alu_shr[23] ;
 wire \alu_shr[24] ;
 wire \alu_shr[25] ;
 wire \alu_shr[26] ;
 wire \alu_shr[27] ;
 wire \alu_shr[28] ;
 wire \alu_shr[29] ;
 wire \alu_shr[2] ;
 wire \alu_shr[30] ;
 wire \alu_shr[31] ;
 wire \alu_shr[3] ;
 wire \alu_shr[4] ;
 wire \alu_shr[5] ;
 wire \alu_shr[6] ;
 wire \alu_shr[7] ;
 wire \alu_shr[8] ;
 wire \alu_shr[9] ;
 wire alu_wait;
 wire \count_cycle[0] ;
 wire \count_cycle[10] ;
 wire \count_cycle[11] ;
 wire \count_cycle[12] ;
 wire \count_cycle[13] ;
 wire \count_cycle[14] ;
 wire \count_cycle[15] ;
 wire \count_cycle[16] ;
 wire \count_cycle[17] ;
 wire \count_cycle[18] ;
 wire \count_cycle[19] ;
 wire \count_cycle[1] ;
 wire \count_cycle[20] ;
 wire \count_cycle[21] ;
 wire \count_cycle[22] ;
 wire \count_cycle[23] ;
 wire \count_cycle[24] ;
 wire \count_cycle[25] ;
 wire \count_cycle[26] ;
 wire \count_cycle[27] ;
 wire \count_cycle[28] ;
 wire \count_cycle[29] ;
 wire \count_cycle[2] ;
 wire \count_cycle[30] ;
 wire \count_cycle[31] ;
 wire \count_cycle[32] ;
 wire \count_cycle[33] ;
 wire \count_cycle[34] ;
 wire \count_cycle[35] ;
 wire \count_cycle[36] ;
 wire \count_cycle[37] ;
 wire \count_cycle[38] ;
 wire \count_cycle[39] ;
 wire \count_cycle[3] ;
 wire \count_cycle[40] ;
 wire \count_cycle[41] ;
 wire \count_cycle[42] ;
 wire \count_cycle[43] ;
 wire \count_cycle[44] ;
 wire \count_cycle[45] ;
 wire \count_cycle[46] ;
 wire \count_cycle[47] ;
 wire \count_cycle[48] ;
 wire \count_cycle[49] ;
 wire \count_cycle[4] ;
 wire \count_cycle[50] ;
 wire \count_cycle[51] ;
 wire \count_cycle[52] ;
 wire \count_cycle[53] ;
 wire \count_cycle[54] ;
 wire \count_cycle[55] ;
 wire \count_cycle[56] ;
 wire \count_cycle[57] ;
 wire \count_cycle[58] ;
 wire \count_cycle[59] ;
 wire \count_cycle[5] ;
 wire \count_cycle[60] ;
 wire \count_cycle[61] ;
 wire \count_cycle[62] ;
 wire \count_cycle[63] ;
 wire \count_cycle[6] ;
 wire \count_cycle[7] ;
 wire \count_cycle[8] ;
 wire \count_cycle[9] ;
 wire \count_instr[0] ;
 wire \count_instr[10] ;
 wire \count_instr[11] ;
 wire \count_instr[12] ;
 wire \count_instr[13] ;
 wire \count_instr[14] ;
 wire \count_instr[15] ;
 wire \count_instr[16] ;
 wire \count_instr[17] ;
 wire \count_instr[18] ;
 wire \count_instr[19] ;
 wire \count_instr[1] ;
 wire \count_instr[20] ;
 wire \count_instr[21] ;
 wire \count_instr[22] ;
 wire \count_instr[23] ;
 wire \count_instr[24] ;
 wire \count_instr[25] ;
 wire \count_instr[26] ;
 wire \count_instr[27] ;
 wire \count_instr[28] ;
 wire \count_instr[29] ;
 wire \count_instr[2] ;
 wire \count_instr[30] ;
 wire \count_instr[31] ;
 wire \count_instr[32] ;
 wire \count_instr[33] ;
 wire \count_instr[34] ;
 wire \count_instr[35] ;
 wire \count_instr[36] ;
 wire \count_instr[37] ;
 wire \count_instr[38] ;
 wire \count_instr[39] ;
 wire \count_instr[3] ;
 wire \count_instr[40] ;
 wire \count_instr[41] ;
 wire \count_instr[42] ;
 wire \count_instr[43] ;
 wire \count_instr[44] ;
 wire \count_instr[45] ;
 wire \count_instr[46] ;
 wire \count_instr[47] ;
 wire \count_instr[48] ;
 wire \count_instr[49] ;
 wire \count_instr[4] ;
 wire \count_instr[50] ;
 wire \count_instr[51] ;
 wire \count_instr[52] ;
 wire \count_instr[53] ;
 wire \count_instr[54] ;
 wire \count_instr[55] ;
 wire \count_instr[56] ;
 wire \count_instr[57] ;
 wire \count_instr[58] ;
 wire \count_instr[59] ;
 wire \count_instr[5] ;
 wire \count_instr[60] ;
 wire \count_instr[61] ;
 wire \count_instr[62] ;
 wire \count_instr[63] ;
 wire \count_instr[6] ;
 wire \count_instr[7] ;
 wire \count_instr[8] ;
 wire \count_instr[9] ;
 wire \cpu_state[0] ;
 wire \cpu_state[1] ;
 wire \cpu_state[2] ;
 wire \cpu_state[3] ;
 wire \cpu_state[4] ;
 wire \cpu_state[5] ;
 wire \cpu_state[6] ;
 wire \cpuregs[0][0] ;
 wire \cpuregs[0][10] ;
 wire \cpuregs[0][11] ;
 wire \cpuregs[0][12] ;
 wire \cpuregs[0][13] ;
 wire \cpuregs[0][14] ;
 wire \cpuregs[0][15] ;
 wire \cpuregs[0][16] ;
 wire \cpuregs[0][17] ;
 wire \cpuregs[0][18] ;
 wire \cpuregs[0][19] ;
 wire \cpuregs[0][1] ;
 wire \cpuregs[0][20] ;
 wire \cpuregs[0][21] ;
 wire \cpuregs[0][22] ;
 wire \cpuregs[0][23] ;
 wire \cpuregs[0][24] ;
 wire \cpuregs[0][25] ;
 wire \cpuregs[0][26] ;
 wire \cpuregs[0][27] ;
 wire \cpuregs[0][28] ;
 wire \cpuregs[0][29] ;
 wire \cpuregs[0][2] ;
 wire \cpuregs[0][30] ;
 wire \cpuregs[0][31] ;
 wire \cpuregs[0][3] ;
 wire \cpuregs[0][4] ;
 wire \cpuregs[0][5] ;
 wire \cpuregs[0][6] ;
 wire \cpuregs[0][7] ;
 wire \cpuregs[0][8] ;
 wire \cpuregs[0][9] ;
 wire \cpuregs[10][0] ;
 wire \cpuregs[10][10] ;
 wire \cpuregs[10][11] ;
 wire \cpuregs[10][12] ;
 wire \cpuregs[10][13] ;
 wire \cpuregs[10][14] ;
 wire \cpuregs[10][15] ;
 wire \cpuregs[10][16] ;
 wire \cpuregs[10][17] ;
 wire \cpuregs[10][18] ;
 wire \cpuregs[10][19] ;
 wire \cpuregs[10][1] ;
 wire \cpuregs[10][20] ;
 wire \cpuregs[10][21] ;
 wire \cpuregs[10][22] ;
 wire \cpuregs[10][23] ;
 wire \cpuregs[10][24] ;
 wire \cpuregs[10][25] ;
 wire \cpuregs[10][26] ;
 wire \cpuregs[10][27] ;
 wire \cpuregs[10][28] ;
 wire \cpuregs[10][29] ;
 wire \cpuregs[10][2] ;
 wire \cpuregs[10][30] ;
 wire \cpuregs[10][31] ;
 wire \cpuregs[10][3] ;
 wire \cpuregs[10][4] ;
 wire \cpuregs[10][5] ;
 wire \cpuregs[10][6] ;
 wire \cpuregs[10][7] ;
 wire \cpuregs[10][8] ;
 wire \cpuregs[10][9] ;
 wire \cpuregs[11][0] ;
 wire \cpuregs[11][10] ;
 wire \cpuregs[11][11] ;
 wire \cpuregs[11][12] ;
 wire \cpuregs[11][13] ;
 wire \cpuregs[11][14] ;
 wire \cpuregs[11][15] ;
 wire \cpuregs[11][16] ;
 wire \cpuregs[11][17] ;
 wire \cpuregs[11][18] ;
 wire \cpuregs[11][19] ;
 wire \cpuregs[11][1] ;
 wire \cpuregs[11][20] ;
 wire \cpuregs[11][21] ;
 wire \cpuregs[11][22] ;
 wire \cpuregs[11][23] ;
 wire \cpuregs[11][24] ;
 wire \cpuregs[11][25] ;
 wire \cpuregs[11][26] ;
 wire \cpuregs[11][27] ;
 wire \cpuregs[11][28] ;
 wire \cpuregs[11][29] ;
 wire \cpuregs[11][2] ;
 wire \cpuregs[11][30] ;
 wire \cpuregs[11][31] ;
 wire \cpuregs[11][3] ;
 wire \cpuregs[11][4] ;
 wire \cpuregs[11][5] ;
 wire \cpuregs[11][6] ;
 wire \cpuregs[11][7] ;
 wire \cpuregs[11][8] ;
 wire \cpuregs[11][9] ;
 wire \cpuregs[12][0] ;
 wire \cpuregs[12][10] ;
 wire \cpuregs[12][11] ;
 wire \cpuregs[12][12] ;
 wire \cpuregs[12][13] ;
 wire \cpuregs[12][14] ;
 wire \cpuregs[12][15] ;
 wire \cpuregs[12][16] ;
 wire \cpuregs[12][17] ;
 wire \cpuregs[12][18] ;
 wire \cpuregs[12][19] ;
 wire \cpuregs[12][1] ;
 wire \cpuregs[12][20] ;
 wire \cpuregs[12][21] ;
 wire \cpuregs[12][22] ;
 wire \cpuregs[12][23] ;
 wire \cpuregs[12][24] ;
 wire \cpuregs[12][25] ;
 wire \cpuregs[12][26] ;
 wire \cpuregs[12][27] ;
 wire \cpuregs[12][28] ;
 wire \cpuregs[12][29] ;
 wire \cpuregs[12][2] ;
 wire \cpuregs[12][30] ;
 wire \cpuregs[12][31] ;
 wire \cpuregs[12][3] ;
 wire \cpuregs[12][4] ;
 wire \cpuregs[12][5] ;
 wire \cpuregs[12][6] ;
 wire \cpuregs[12][7] ;
 wire \cpuregs[12][8] ;
 wire \cpuregs[12][9] ;
 wire \cpuregs[13][0] ;
 wire \cpuregs[13][10] ;
 wire \cpuregs[13][11] ;
 wire \cpuregs[13][12] ;
 wire \cpuregs[13][13] ;
 wire \cpuregs[13][14] ;
 wire \cpuregs[13][15] ;
 wire \cpuregs[13][16] ;
 wire \cpuregs[13][17] ;
 wire \cpuregs[13][18] ;
 wire \cpuregs[13][19] ;
 wire \cpuregs[13][1] ;
 wire \cpuregs[13][20] ;
 wire \cpuregs[13][21] ;
 wire \cpuregs[13][22] ;
 wire \cpuregs[13][23] ;
 wire \cpuregs[13][24] ;
 wire \cpuregs[13][25] ;
 wire \cpuregs[13][26] ;
 wire \cpuregs[13][27] ;
 wire \cpuregs[13][28] ;
 wire \cpuregs[13][29] ;
 wire \cpuregs[13][2] ;
 wire \cpuregs[13][30] ;
 wire \cpuregs[13][31] ;
 wire \cpuregs[13][3] ;
 wire \cpuregs[13][4] ;
 wire \cpuregs[13][5] ;
 wire \cpuregs[13][6] ;
 wire \cpuregs[13][7] ;
 wire \cpuregs[13][8] ;
 wire \cpuregs[13][9] ;
 wire \cpuregs[14][0] ;
 wire \cpuregs[14][10] ;
 wire \cpuregs[14][11] ;
 wire \cpuregs[14][12] ;
 wire \cpuregs[14][13] ;
 wire \cpuregs[14][14] ;
 wire \cpuregs[14][15] ;
 wire \cpuregs[14][16] ;
 wire \cpuregs[14][17] ;
 wire \cpuregs[14][18] ;
 wire \cpuregs[14][19] ;
 wire \cpuregs[14][1] ;
 wire \cpuregs[14][20] ;
 wire \cpuregs[14][21] ;
 wire \cpuregs[14][22] ;
 wire \cpuregs[14][23] ;
 wire \cpuregs[14][24] ;
 wire \cpuregs[14][25] ;
 wire \cpuregs[14][26] ;
 wire \cpuregs[14][27] ;
 wire \cpuregs[14][28] ;
 wire \cpuregs[14][29] ;
 wire \cpuregs[14][2] ;
 wire \cpuregs[14][30] ;
 wire \cpuregs[14][31] ;
 wire \cpuregs[14][3] ;
 wire \cpuregs[14][4] ;
 wire \cpuregs[14][5] ;
 wire \cpuregs[14][6] ;
 wire \cpuregs[14][7] ;
 wire \cpuregs[14][8] ;
 wire \cpuregs[14][9] ;
 wire \cpuregs[15][0] ;
 wire \cpuregs[15][10] ;
 wire \cpuregs[15][11] ;
 wire \cpuregs[15][12] ;
 wire \cpuregs[15][13] ;
 wire \cpuregs[15][14] ;
 wire \cpuregs[15][15] ;
 wire \cpuregs[15][16] ;
 wire \cpuregs[15][17] ;
 wire \cpuregs[15][18] ;
 wire \cpuregs[15][19] ;
 wire \cpuregs[15][1] ;
 wire \cpuregs[15][20] ;
 wire \cpuregs[15][21] ;
 wire \cpuregs[15][22] ;
 wire \cpuregs[15][23] ;
 wire \cpuregs[15][24] ;
 wire \cpuregs[15][25] ;
 wire \cpuregs[15][26] ;
 wire \cpuregs[15][27] ;
 wire \cpuregs[15][28] ;
 wire \cpuregs[15][29] ;
 wire \cpuregs[15][2] ;
 wire \cpuregs[15][30] ;
 wire \cpuregs[15][31] ;
 wire \cpuregs[15][3] ;
 wire \cpuregs[15][4] ;
 wire \cpuregs[15][5] ;
 wire \cpuregs[15][6] ;
 wire \cpuregs[15][7] ;
 wire \cpuregs[15][8] ;
 wire \cpuregs[15][9] ;
 wire \cpuregs[16][0] ;
 wire \cpuregs[16][10] ;
 wire \cpuregs[16][11] ;
 wire \cpuregs[16][12] ;
 wire \cpuregs[16][13] ;
 wire \cpuregs[16][14] ;
 wire \cpuregs[16][15] ;
 wire \cpuregs[16][16] ;
 wire \cpuregs[16][17] ;
 wire \cpuregs[16][18] ;
 wire \cpuregs[16][19] ;
 wire \cpuregs[16][1] ;
 wire \cpuregs[16][20] ;
 wire \cpuregs[16][21] ;
 wire \cpuregs[16][22] ;
 wire \cpuregs[16][23] ;
 wire \cpuregs[16][24] ;
 wire \cpuregs[16][25] ;
 wire \cpuregs[16][26] ;
 wire \cpuregs[16][27] ;
 wire \cpuregs[16][28] ;
 wire \cpuregs[16][29] ;
 wire \cpuregs[16][2] ;
 wire \cpuregs[16][30] ;
 wire \cpuregs[16][31] ;
 wire \cpuregs[16][3] ;
 wire \cpuregs[16][4] ;
 wire \cpuregs[16][5] ;
 wire \cpuregs[16][6] ;
 wire \cpuregs[16][7] ;
 wire \cpuregs[16][8] ;
 wire \cpuregs[16][9] ;
 wire \cpuregs[17][0] ;
 wire \cpuregs[17][10] ;
 wire \cpuregs[17][11] ;
 wire \cpuregs[17][12] ;
 wire \cpuregs[17][13] ;
 wire \cpuregs[17][14] ;
 wire \cpuregs[17][15] ;
 wire \cpuregs[17][16] ;
 wire \cpuregs[17][17] ;
 wire \cpuregs[17][18] ;
 wire \cpuregs[17][19] ;
 wire \cpuregs[17][1] ;
 wire \cpuregs[17][20] ;
 wire \cpuregs[17][21] ;
 wire \cpuregs[17][22] ;
 wire \cpuregs[17][23] ;
 wire \cpuregs[17][24] ;
 wire \cpuregs[17][25] ;
 wire \cpuregs[17][26] ;
 wire \cpuregs[17][27] ;
 wire \cpuregs[17][28] ;
 wire \cpuregs[17][29] ;
 wire \cpuregs[17][2] ;
 wire \cpuregs[17][30] ;
 wire \cpuregs[17][31] ;
 wire \cpuregs[17][3] ;
 wire \cpuregs[17][4] ;
 wire \cpuregs[17][5] ;
 wire \cpuregs[17][6] ;
 wire \cpuregs[17][7] ;
 wire \cpuregs[17][8] ;
 wire \cpuregs[17][9] ;
 wire \cpuregs[18][0] ;
 wire \cpuregs[18][10] ;
 wire \cpuregs[18][11] ;
 wire \cpuregs[18][12] ;
 wire \cpuregs[18][13] ;
 wire \cpuregs[18][14] ;
 wire \cpuregs[18][15] ;
 wire \cpuregs[18][16] ;
 wire \cpuregs[18][17] ;
 wire \cpuregs[18][18] ;
 wire \cpuregs[18][19] ;
 wire \cpuregs[18][1] ;
 wire \cpuregs[18][20] ;
 wire \cpuregs[18][21] ;
 wire \cpuregs[18][22] ;
 wire \cpuregs[18][23] ;
 wire \cpuregs[18][24] ;
 wire \cpuregs[18][25] ;
 wire \cpuregs[18][26] ;
 wire \cpuregs[18][27] ;
 wire \cpuregs[18][28] ;
 wire \cpuregs[18][29] ;
 wire \cpuregs[18][2] ;
 wire \cpuregs[18][30] ;
 wire \cpuregs[18][31] ;
 wire \cpuregs[18][3] ;
 wire \cpuregs[18][4] ;
 wire \cpuregs[18][5] ;
 wire \cpuregs[18][6] ;
 wire \cpuregs[18][7] ;
 wire \cpuregs[18][8] ;
 wire \cpuregs[18][9] ;
 wire \cpuregs[19][0] ;
 wire \cpuregs[19][10] ;
 wire \cpuregs[19][11] ;
 wire \cpuregs[19][12] ;
 wire \cpuregs[19][13] ;
 wire \cpuregs[19][14] ;
 wire \cpuregs[19][15] ;
 wire \cpuregs[19][16] ;
 wire \cpuregs[19][17] ;
 wire \cpuregs[19][18] ;
 wire \cpuregs[19][19] ;
 wire \cpuregs[19][1] ;
 wire \cpuregs[19][20] ;
 wire \cpuregs[19][21] ;
 wire \cpuregs[19][22] ;
 wire \cpuregs[19][23] ;
 wire \cpuregs[19][24] ;
 wire \cpuregs[19][25] ;
 wire \cpuregs[19][26] ;
 wire \cpuregs[19][27] ;
 wire \cpuregs[19][28] ;
 wire \cpuregs[19][29] ;
 wire \cpuregs[19][2] ;
 wire \cpuregs[19][30] ;
 wire \cpuregs[19][31] ;
 wire \cpuregs[19][3] ;
 wire \cpuregs[19][4] ;
 wire \cpuregs[19][5] ;
 wire \cpuregs[19][6] ;
 wire \cpuregs[19][7] ;
 wire \cpuregs[19][8] ;
 wire \cpuregs[19][9] ;
 wire \cpuregs[1][0] ;
 wire \cpuregs[1][10] ;
 wire \cpuregs[1][11] ;
 wire \cpuregs[1][12] ;
 wire \cpuregs[1][13] ;
 wire \cpuregs[1][14] ;
 wire \cpuregs[1][15] ;
 wire \cpuregs[1][16] ;
 wire \cpuregs[1][17] ;
 wire \cpuregs[1][18] ;
 wire \cpuregs[1][19] ;
 wire \cpuregs[1][1] ;
 wire \cpuregs[1][20] ;
 wire \cpuregs[1][21] ;
 wire \cpuregs[1][22] ;
 wire \cpuregs[1][23] ;
 wire \cpuregs[1][24] ;
 wire \cpuregs[1][25] ;
 wire \cpuregs[1][26] ;
 wire \cpuregs[1][27] ;
 wire \cpuregs[1][28] ;
 wire \cpuregs[1][29] ;
 wire \cpuregs[1][2] ;
 wire \cpuregs[1][30] ;
 wire \cpuregs[1][31] ;
 wire \cpuregs[1][3] ;
 wire \cpuregs[1][4] ;
 wire \cpuregs[1][5] ;
 wire \cpuregs[1][6] ;
 wire \cpuregs[1][7] ;
 wire \cpuregs[1][8] ;
 wire \cpuregs[1][9] ;
 wire \cpuregs[2][0] ;
 wire \cpuregs[2][10] ;
 wire \cpuregs[2][11] ;
 wire \cpuregs[2][12] ;
 wire \cpuregs[2][13] ;
 wire \cpuregs[2][14] ;
 wire \cpuregs[2][15] ;
 wire \cpuregs[2][16] ;
 wire \cpuregs[2][17] ;
 wire \cpuregs[2][18] ;
 wire \cpuregs[2][19] ;
 wire \cpuregs[2][1] ;
 wire \cpuregs[2][20] ;
 wire \cpuregs[2][21] ;
 wire \cpuregs[2][22] ;
 wire \cpuregs[2][23] ;
 wire \cpuregs[2][24] ;
 wire \cpuregs[2][25] ;
 wire \cpuregs[2][26] ;
 wire \cpuregs[2][27] ;
 wire \cpuregs[2][28] ;
 wire \cpuregs[2][29] ;
 wire \cpuregs[2][2] ;
 wire \cpuregs[2][30] ;
 wire \cpuregs[2][31] ;
 wire \cpuregs[2][3] ;
 wire \cpuregs[2][4] ;
 wire \cpuregs[2][5] ;
 wire \cpuregs[2][6] ;
 wire \cpuregs[2][7] ;
 wire \cpuregs[2][8] ;
 wire \cpuregs[2][9] ;
 wire \cpuregs[3][0] ;
 wire \cpuregs[3][10] ;
 wire \cpuregs[3][11] ;
 wire \cpuregs[3][12] ;
 wire \cpuregs[3][13] ;
 wire \cpuregs[3][14] ;
 wire \cpuregs[3][15] ;
 wire \cpuregs[3][16] ;
 wire \cpuregs[3][17] ;
 wire \cpuregs[3][18] ;
 wire \cpuregs[3][19] ;
 wire \cpuregs[3][1] ;
 wire \cpuregs[3][20] ;
 wire \cpuregs[3][21] ;
 wire \cpuregs[3][22] ;
 wire \cpuregs[3][23] ;
 wire \cpuregs[3][24] ;
 wire \cpuregs[3][25] ;
 wire \cpuregs[3][26] ;
 wire \cpuregs[3][27] ;
 wire \cpuregs[3][28] ;
 wire \cpuregs[3][29] ;
 wire \cpuregs[3][2] ;
 wire \cpuregs[3][30] ;
 wire \cpuregs[3][31] ;
 wire \cpuregs[3][3] ;
 wire \cpuregs[3][4] ;
 wire \cpuregs[3][5] ;
 wire \cpuregs[3][6] ;
 wire \cpuregs[3][7] ;
 wire \cpuregs[3][8] ;
 wire \cpuregs[3][9] ;
 wire \cpuregs[4][0] ;
 wire \cpuregs[4][10] ;
 wire \cpuregs[4][11] ;
 wire \cpuregs[4][12] ;
 wire \cpuregs[4][13] ;
 wire \cpuregs[4][14] ;
 wire \cpuregs[4][15] ;
 wire \cpuregs[4][16] ;
 wire \cpuregs[4][17] ;
 wire \cpuregs[4][18] ;
 wire \cpuregs[4][19] ;
 wire \cpuregs[4][1] ;
 wire \cpuregs[4][20] ;
 wire \cpuregs[4][21] ;
 wire \cpuregs[4][22] ;
 wire \cpuregs[4][23] ;
 wire \cpuregs[4][24] ;
 wire \cpuregs[4][25] ;
 wire \cpuregs[4][26] ;
 wire \cpuregs[4][27] ;
 wire \cpuregs[4][28] ;
 wire \cpuregs[4][29] ;
 wire \cpuregs[4][2] ;
 wire \cpuregs[4][30] ;
 wire \cpuregs[4][31] ;
 wire \cpuregs[4][3] ;
 wire \cpuregs[4][4] ;
 wire \cpuregs[4][5] ;
 wire \cpuregs[4][6] ;
 wire \cpuregs[4][7] ;
 wire \cpuregs[4][8] ;
 wire \cpuregs[4][9] ;
 wire \cpuregs[5][0] ;
 wire \cpuregs[5][10] ;
 wire \cpuregs[5][11] ;
 wire \cpuregs[5][12] ;
 wire \cpuregs[5][13] ;
 wire \cpuregs[5][14] ;
 wire \cpuregs[5][15] ;
 wire \cpuregs[5][16] ;
 wire \cpuregs[5][17] ;
 wire \cpuregs[5][18] ;
 wire \cpuregs[5][19] ;
 wire \cpuregs[5][1] ;
 wire \cpuregs[5][20] ;
 wire \cpuregs[5][21] ;
 wire \cpuregs[5][22] ;
 wire \cpuregs[5][23] ;
 wire \cpuregs[5][24] ;
 wire \cpuregs[5][25] ;
 wire \cpuregs[5][26] ;
 wire \cpuregs[5][27] ;
 wire \cpuregs[5][28] ;
 wire \cpuregs[5][29] ;
 wire \cpuregs[5][2] ;
 wire \cpuregs[5][30] ;
 wire \cpuregs[5][31] ;
 wire \cpuregs[5][3] ;
 wire \cpuregs[5][4] ;
 wire \cpuregs[5][5] ;
 wire \cpuregs[5][6] ;
 wire \cpuregs[5][7] ;
 wire \cpuregs[5][8] ;
 wire \cpuregs[5][9] ;
 wire \cpuregs[6][0] ;
 wire \cpuregs[6][10] ;
 wire \cpuregs[6][11] ;
 wire \cpuregs[6][12] ;
 wire \cpuregs[6][13] ;
 wire \cpuregs[6][14] ;
 wire \cpuregs[6][15] ;
 wire \cpuregs[6][16] ;
 wire \cpuregs[6][17] ;
 wire \cpuregs[6][18] ;
 wire \cpuregs[6][19] ;
 wire \cpuregs[6][1] ;
 wire \cpuregs[6][20] ;
 wire \cpuregs[6][21] ;
 wire \cpuregs[6][22] ;
 wire \cpuregs[6][23] ;
 wire \cpuregs[6][24] ;
 wire \cpuregs[6][25] ;
 wire \cpuregs[6][26] ;
 wire \cpuregs[6][27] ;
 wire \cpuregs[6][28] ;
 wire \cpuregs[6][29] ;
 wire \cpuregs[6][2] ;
 wire \cpuregs[6][30] ;
 wire \cpuregs[6][31] ;
 wire \cpuregs[6][3] ;
 wire \cpuregs[6][4] ;
 wire \cpuregs[6][5] ;
 wire \cpuregs[6][6] ;
 wire \cpuregs[6][7] ;
 wire \cpuregs[6][8] ;
 wire \cpuregs[6][9] ;
 wire \cpuregs[7][0] ;
 wire \cpuregs[7][10] ;
 wire \cpuregs[7][11] ;
 wire \cpuregs[7][12] ;
 wire \cpuregs[7][13] ;
 wire \cpuregs[7][14] ;
 wire \cpuregs[7][15] ;
 wire \cpuregs[7][16] ;
 wire \cpuregs[7][17] ;
 wire \cpuregs[7][18] ;
 wire \cpuregs[7][19] ;
 wire \cpuregs[7][1] ;
 wire \cpuregs[7][20] ;
 wire \cpuregs[7][21] ;
 wire \cpuregs[7][22] ;
 wire \cpuregs[7][23] ;
 wire \cpuregs[7][24] ;
 wire \cpuregs[7][25] ;
 wire \cpuregs[7][26] ;
 wire \cpuregs[7][27] ;
 wire \cpuregs[7][28] ;
 wire \cpuregs[7][29] ;
 wire \cpuregs[7][2] ;
 wire \cpuregs[7][30] ;
 wire \cpuregs[7][31] ;
 wire \cpuregs[7][3] ;
 wire \cpuregs[7][4] ;
 wire \cpuregs[7][5] ;
 wire \cpuregs[7][6] ;
 wire \cpuregs[7][7] ;
 wire \cpuregs[7][8] ;
 wire \cpuregs[7][9] ;
 wire \cpuregs[8][0] ;
 wire \cpuregs[8][10] ;
 wire \cpuregs[8][11] ;
 wire \cpuregs[8][12] ;
 wire \cpuregs[8][13] ;
 wire \cpuregs[8][14] ;
 wire \cpuregs[8][15] ;
 wire \cpuregs[8][16] ;
 wire \cpuregs[8][17] ;
 wire \cpuregs[8][18] ;
 wire \cpuregs[8][19] ;
 wire \cpuregs[8][1] ;
 wire \cpuregs[8][20] ;
 wire \cpuregs[8][21] ;
 wire \cpuregs[8][22] ;
 wire \cpuregs[8][23] ;
 wire \cpuregs[8][24] ;
 wire \cpuregs[8][25] ;
 wire \cpuregs[8][26] ;
 wire \cpuregs[8][27] ;
 wire \cpuregs[8][28] ;
 wire \cpuregs[8][29] ;
 wire \cpuregs[8][2] ;
 wire \cpuregs[8][30] ;
 wire \cpuregs[8][31] ;
 wire \cpuregs[8][3] ;
 wire \cpuregs[8][4] ;
 wire \cpuregs[8][5] ;
 wire \cpuregs[8][6] ;
 wire \cpuregs[8][7] ;
 wire \cpuregs[8][8] ;
 wire \cpuregs[8][9] ;
 wire \cpuregs[9][0] ;
 wire \cpuregs[9][10] ;
 wire \cpuregs[9][11] ;
 wire \cpuregs[9][12] ;
 wire \cpuregs[9][13] ;
 wire \cpuregs[9][14] ;
 wire \cpuregs[9][15] ;
 wire \cpuregs[9][16] ;
 wire \cpuregs[9][17] ;
 wire \cpuregs[9][18] ;
 wire \cpuregs[9][19] ;
 wire \cpuregs[9][1] ;
 wire \cpuregs[9][20] ;
 wire \cpuregs[9][21] ;
 wire \cpuregs[9][22] ;
 wire \cpuregs[9][23] ;
 wire \cpuregs[9][24] ;
 wire \cpuregs[9][25] ;
 wire \cpuregs[9][26] ;
 wire \cpuregs[9][27] ;
 wire \cpuregs[9][28] ;
 wire \cpuregs[9][29] ;
 wire \cpuregs[9][2] ;
 wire \cpuregs[9][30] ;
 wire \cpuregs[9][31] ;
 wire \cpuregs[9][3] ;
 wire \cpuregs[9][4] ;
 wire \cpuregs[9][5] ;
 wire \cpuregs[9][6] ;
 wire \cpuregs[9][7] ;
 wire \cpuregs[9][8] ;
 wire \cpuregs[9][9] ;
 wire \decoded_imm[0] ;
 wire \decoded_imm[10] ;
 wire \decoded_imm[11] ;
 wire \decoded_imm[12] ;
 wire \decoded_imm[13] ;
 wire \decoded_imm[14] ;
 wire \decoded_imm[15] ;
 wire \decoded_imm[16] ;
 wire \decoded_imm[17] ;
 wire \decoded_imm[18] ;
 wire \decoded_imm[19] ;
 wire \decoded_imm[1] ;
 wire \decoded_imm[20] ;
 wire \decoded_imm[21] ;
 wire \decoded_imm[22] ;
 wire \decoded_imm[23] ;
 wire \decoded_imm[24] ;
 wire \decoded_imm[25] ;
 wire \decoded_imm[26] ;
 wire \decoded_imm[27] ;
 wire \decoded_imm[28] ;
 wire \decoded_imm[29] ;
 wire \decoded_imm[2] ;
 wire \decoded_imm[30] ;
 wire \decoded_imm[31] ;
 wire \decoded_imm[3] ;
 wire \decoded_imm[4] ;
 wire \decoded_imm[5] ;
 wire \decoded_imm[6] ;
 wire \decoded_imm[7] ;
 wire \decoded_imm[8] ;
 wire \decoded_imm[9] ;
 wire \decoded_imm_uj[10] ;
 wire \decoded_imm_uj[11] ;
 wire \decoded_imm_uj[12] ;
 wire \decoded_imm_uj[13] ;
 wire \decoded_imm_uj[14] ;
 wire \decoded_imm_uj[15] ;
 wire \decoded_imm_uj[16] ;
 wire \decoded_imm_uj[17] ;
 wire \decoded_imm_uj[18] ;
 wire \decoded_imm_uj[19] ;
 wire \decoded_imm_uj[1] ;
 wire \decoded_imm_uj[20] ;
 wire \decoded_imm_uj[2] ;
 wire \decoded_imm_uj[3] ;
 wire \decoded_imm_uj[4] ;
 wire \decoded_imm_uj[5] ;
 wire \decoded_imm_uj[6] ;
 wire \decoded_imm_uj[7] ;
 wire \decoded_imm_uj[8] ;
 wire \decoded_imm_uj[9] ;
 wire \decoded_rd[0] ;
 wire \decoded_rd[1] ;
 wire \decoded_rd[2] ;
 wire \decoded_rd[3] ;
 wire \decoded_rd[4] ;
 wire \decoded_rs1[0] ;
 wire \decoded_rs1[1] ;
 wire \decoded_rs1[2] ;
 wire \decoded_rs1[3] ;
 wire \decoded_rs1[4] ;
 wire decoder_pseudo_trigger;
 wire decoder_trigger;
 wire do_waitirq;
 wire \genblk1.pcpi_mul.active[0] ;
 wire \genblk1.pcpi_mul.active[1] ;
 wire \genblk1.pcpi_mul.instr_any_mulh ;
 wire \genblk1.pcpi_mul.rd[0] ;
 wire \genblk1.pcpi_mul.rd[10] ;
 wire \genblk1.pcpi_mul.rd[11] ;
 wire \genblk1.pcpi_mul.rd[12] ;
 wire \genblk1.pcpi_mul.rd[13] ;
 wire \genblk1.pcpi_mul.rd[14] ;
 wire \genblk1.pcpi_mul.rd[15] ;
 wire \genblk1.pcpi_mul.rd[16] ;
 wire \genblk1.pcpi_mul.rd[17] ;
 wire \genblk1.pcpi_mul.rd[18] ;
 wire \genblk1.pcpi_mul.rd[19] ;
 wire \genblk1.pcpi_mul.rd[1] ;
 wire \genblk1.pcpi_mul.rd[20] ;
 wire \genblk1.pcpi_mul.rd[21] ;
 wire \genblk1.pcpi_mul.rd[22] ;
 wire \genblk1.pcpi_mul.rd[23] ;
 wire \genblk1.pcpi_mul.rd[24] ;
 wire \genblk1.pcpi_mul.rd[25] ;
 wire \genblk1.pcpi_mul.rd[26] ;
 wire \genblk1.pcpi_mul.rd[27] ;
 wire \genblk1.pcpi_mul.rd[28] ;
 wire \genblk1.pcpi_mul.rd[29] ;
 wire \genblk1.pcpi_mul.rd[2] ;
 wire \genblk1.pcpi_mul.rd[30] ;
 wire \genblk1.pcpi_mul.rd[31] ;
 wire \genblk1.pcpi_mul.rd[32] ;
 wire \genblk1.pcpi_mul.rd[33] ;
 wire \genblk1.pcpi_mul.rd[34] ;
 wire \genblk1.pcpi_mul.rd[35] ;
 wire \genblk1.pcpi_mul.rd[36] ;
 wire \genblk1.pcpi_mul.rd[37] ;
 wire \genblk1.pcpi_mul.rd[38] ;
 wire \genblk1.pcpi_mul.rd[39] ;
 wire \genblk1.pcpi_mul.rd[3] ;
 wire \genblk1.pcpi_mul.rd[40] ;
 wire \genblk1.pcpi_mul.rd[41] ;
 wire \genblk1.pcpi_mul.rd[42] ;
 wire \genblk1.pcpi_mul.rd[43] ;
 wire \genblk1.pcpi_mul.rd[44] ;
 wire \genblk1.pcpi_mul.rd[45] ;
 wire \genblk1.pcpi_mul.rd[46] ;
 wire \genblk1.pcpi_mul.rd[47] ;
 wire \genblk1.pcpi_mul.rd[48] ;
 wire \genblk1.pcpi_mul.rd[49] ;
 wire \genblk1.pcpi_mul.rd[4] ;
 wire \genblk1.pcpi_mul.rd[50] ;
 wire \genblk1.pcpi_mul.rd[51] ;
 wire \genblk1.pcpi_mul.rd[52] ;
 wire \genblk1.pcpi_mul.rd[53] ;
 wire \genblk1.pcpi_mul.rd[54] ;
 wire \genblk1.pcpi_mul.rd[55] ;
 wire \genblk1.pcpi_mul.rd[56] ;
 wire \genblk1.pcpi_mul.rd[57] ;
 wire \genblk1.pcpi_mul.rd[58] ;
 wire \genblk1.pcpi_mul.rd[59] ;
 wire \genblk1.pcpi_mul.rd[5] ;
 wire \genblk1.pcpi_mul.rd[60] ;
 wire \genblk1.pcpi_mul.rd[61] ;
 wire \genblk1.pcpi_mul.rd[62] ;
 wire \genblk1.pcpi_mul.rd[63] ;
 wire \genblk1.pcpi_mul.rd[6] ;
 wire \genblk1.pcpi_mul.rd[7] ;
 wire \genblk1.pcpi_mul.rd[8] ;
 wire \genblk1.pcpi_mul.rd[9] ;
 wire \genblk1.pcpi_mul.rs1[0] ;
 wire \genblk1.pcpi_mul.rs1[10] ;
 wire \genblk1.pcpi_mul.rs1[11] ;
 wire \genblk1.pcpi_mul.rs1[12] ;
 wire \genblk1.pcpi_mul.rs1[13] ;
 wire \genblk1.pcpi_mul.rs1[14] ;
 wire \genblk1.pcpi_mul.rs1[15] ;
 wire \genblk1.pcpi_mul.rs1[16] ;
 wire \genblk1.pcpi_mul.rs1[17] ;
 wire \genblk1.pcpi_mul.rs1[18] ;
 wire \genblk1.pcpi_mul.rs1[19] ;
 wire \genblk1.pcpi_mul.rs1[1] ;
 wire \genblk1.pcpi_mul.rs1[20] ;
 wire \genblk1.pcpi_mul.rs1[21] ;
 wire \genblk1.pcpi_mul.rs1[22] ;
 wire \genblk1.pcpi_mul.rs1[23] ;
 wire \genblk1.pcpi_mul.rs1[24] ;
 wire \genblk1.pcpi_mul.rs1[25] ;
 wire \genblk1.pcpi_mul.rs1[26] ;
 wire \genblk1.pcpi_mul.rs1[27] ;
 wire \genblk1.pcpi_mul.rs1[28] ;
 wire \genblk1.pcpi_mul.rs1[29] ;
 wire \genblk1.pcpi_mul.rs1[2] ;
 wire \genblk1.pcpi_mul.rs1[30] ;
 wire \genblk1.pcpi_mul.rs1[31] ;
 wire \genblk1.pcpi_mul.rs1[32] ;
 wire \genblk1.pcpi_mul.rs1[3] ;
 wire \genblk1.pcpi_mul.rs1[4] ;
 wire \genblk1.pcpi_mul.rs1[5] ;
 wire \genblk1.pcpi_mul.rs1[6] ;
 wire \genblk1.pcpi_mul.rs1[7] ;
 wire \genblk1.pcpi_mul.rs1[8] ;
 wire \genblk1.pcpi_mul.rs1[9] ;
 wire \genblk1.pcpi_mul.rs2[0] ;
 wire \genblk1.pcpi_mul.rs2[10] ;
 wire \genblk1.pcpi_mul.rs2[11] ;
 wire \genblk1.pcpi_mul.rs2[12] ;
 wire \genblk1.pcpi_mul.rs2[13] ;
 wire \genblk1.pcpi_mul.rs2[14] ;
 wire \genblk1.pcpi_mul.rs2[15] ;
 wire \genblk1.pcpi_mul.rs2[16] ;
 wire \genblk1.pcpi_mul.rs2[17] ;
 wire \genblk1.pcpi_mul.rs2[18] ;
 wire \genblk1.pcpi_mul.rs2[19] ;
 wire \genblk1.pcpi_mul.rs2[1] ;
 wire \genblk1.pcpi_mul.rs2[20] ;
 wire \genblk1.pcpi_mul.rs2[21] ;
 wire \genblk1.pcpi_mul.rs2[22] ;
 wire \genblk1.pcpi_mul.rs2[23] ;
 wire \genblk1.pcpi_mul.rs2[24] ;
 wire \genblk1.pcpi_mul.rs2[25] ;
 wire \genblk1.pcpi_mul.rs2[26] ;
 wire \genblk1.pcpi_mul.rs2[27] ;
 wire \genblk1.pcpi_mul.rs2[28] ;
 wire \genblk1.pcpi_mul.rs2[29] ;
 wire \genblk1.pcpi_mul.rs2[2] ;
 wire \genblk1.pcpi_mul.rs2[30] ;
 wire \genblk1.pcpi_mul.rs2[31] ;
 wire \genblk1.pcpi_mul.rs2[32] ;
 wire \genblk1.pcpi_mul.rs2[3] ;
 wire \genblk1.pcpi_mul.rs2[4] ;
 wire \genblk1.pcpi_mul.rs2[5] ;
 wire \genblk1.pcpi_mul.rs2[6] ;
 wire \genblk1.pcpi_mul.rs2[7] ;
 wire \genblk1.pcpi_mul.rs2[8] ;
 wire \genblk1.pcpi_mul.rs2[9] ;
 wire \genblk1.pcpi_mul.shift_out ;
 wire instr_add;
 wire instr_addi;
 wire instr_and;
 wire instr_andi;
 wire instr_auipc;
 wire instr_beq;
 wire instr_bge;
 wire instr_bgeu;
 wire instr_blt;
 wire instr_bltu;
 wire instr_bne;
 wire instr_ecall_ebreak;
 wire instr_getq;
 wire instr_jal;
 wire instr_jalr;
 wire instr_lb;
 wire instr_lbu;
 wire instr_lh;
 wire instr_lhu;
 wire instr_lui;
 wire instr_lw;
 wire instr_maskirq;
 wire instr_or;
 wire instr_ori;
 wire instr_rdcycle;
 wire instr_rdcycleh;
 wire instr_rdinstr;
 wire instr_rdinstrh;
 wire instr_retirq;
 wire instr_sb;
 wire instr_setq;
 wire instr_sh;
 wire instr_sll;
 wire instr_slli;
 wire instr_slt;
 wire instr_slti;
 wire instr_sltiu;
 wire instr_sltu;
 wire instr_sra;
 wire instr_srai;
 wire instr_srl;
 wire instr_srli;
 wire instr_sub;
 wire instr_sw;
 wire instr_timer;
 wire instr_waitirq;
 wire instr_xor;
 wire instr_xori;
 wire irq_active;
 wire irq_delay;
 wire \irq_mask[0] ;
 wire \irq_mask[10] ;
 wire \irq_mask[11] ;
 wire \irq_mask[12] ;
 wire \irq_mask[13] ;
 wire \irq_mask[14] ;
 wire \irq_mask[15] ;
 wire \irq_mask[16] ;
 wire \irq_mask[17] ;
 wire \irq_mask[18] ;
 wire \irq_mask[19] ;
 wire \irq_mask[1] ;
 wire \irq_mask[20] ;
 wire \irq_mask[21] ;
 wire \irq_mask[22] ;
 wire \irq_mask[23] ;
 wire \irq_mask[24] ;
 wire \irq_mask[25] ;
 wire \irq_mask[26] ;
 wire \irq_mask[27] ;
 wire \irq_mask[28] ;
 wire \irq_mask[29] ;
 wire \irq_mask[2] ;
 wire \irq_mask[30] ;
 wire \irq_mask[31] ;
 wire \irq_mask[3] ;
 wire \irq_mask[4] ;
 wire \irq_mask[5] ;
 wire \irq_mask[6] ;
 wire \irq_mask[7] ;
 wire \irq_mask[8] ;
 wire \irq_mask[9] ;
 wire \irq_pending[0] ;
 wire \irq_pending[10] ;
 wire \irq_pending[11] ;
 wire \irq_pending[12] ;
 wire \irq_pending[13] ;
 wire \irq_pending[14] ;
 wire \irq_pending[15] ;
 wire \irq_pending[16] ;
 wire \irq_pending[17] ;
 wire \irq_pending[18] ;
 wire \irq_pending[19] ;
 wire \irq_pending[1] ;
 wire \irq_pending[20] ;
 wire \irq_pending[21] ;
 wire \irq_pending[22] ;
 wire \irq_pending[23] ;
 wire \irq_pending[24] ;
 wire \irq_pending[25] ;
 wire \irq_pending[26] ;
 wire \irq_pending[27] ;
 wire \irq_pending[28] ;
 wire \irq_pending[29] ;
 wire \irq_pending[2] ;
 wire \irq_pending[30] ;
 wire \irq_pending[31] ;
 wire \irq_pending[3] ;
 wire \irq_pending[4] ;
 wire \irq_pending[5] ;
 wire \irq_pending[6] ;
 wire \irq_pending[7] ;
 wire \irq_pending[8] ;
 wire \irq_pending[9] ;
 wire \irq_state[0] ;
 wire \irq_state[1] ;
 wire is_alu_reg_imm;
 wire is_alu_reg_reg;
 wire is_beq_bne_blt_bge_bltu_bgeu;
 wire is_compare;
 wire is_jalr_addi_slti_sltiu_xori_ori_andi;
 wire is_lb_lh_lw_lbu_lhu;
 wire is_lui_auipc_jal;
 wire is_sb_sh_sw;
 wire is_slli_srli_srai;
 wire is_slti_blt_slt;
 wire is_sltiu_bltu_sltu;
 wire latched_branch;
 wire latched_is_lb;
 wire latched_is_lh;
 wire \latched_rd[0] ;
 wire \latched_rd[1] ;
 wire \latched_rd[2] ;
 wire \latched_rd[3] ;
 wire \latched_rd[4] ;
 wire latched_stalu;
 wire latched_store;
 wire net375;
 wire net376;
 wire mem_do_prefetch;
 wire mem_do_rdata;
 wire mem_do_rinst;
 wire mem_do_wdata;
 wire net377;
 wire net378;
 wire \mem_rdata_q[0] ;
 wire \mem_rdata_q[10] ;
 wire \mem_rdata_q[11] ;
 wire \mem_rdata_q[12] ;
 wire \mem_rdata_q[13] ;
 wire \mem_rdata_q[14] ;
 wire \mem_rdata_q[15] ;
 wire \mem_rdata_q[16] ;
 wire \mem_rdata_q[17] ;
 wire \mem_rdata_q[18] ;
 wire \mem_rdata_q[19] ;
 wire \mem_rdata_q[1] ;
 wire \mem_rdata_q[20] ;
 wire \mem_rdata_q[21] ;
 wire \mem_rdata_q[22] ;
 wire \mem_rdata_q[23] ;
 wire \mem_rdata_q[24] ;
 wire \mem_rdata_q[25] ;
 wire \mem_rdata_q[26] ;
 wire \mem_rdata_q[27] ;
 wire \mem_rdata_q[28] ;
 wire \mem_rdata_q[29] ;
 wire \mem_rdata_q[2] ;
 wire \mem_rdata_q[30] ;
 wire \mem_rdata_q[31] ;
 wire \mem_rdata_q[3] ;
 wire \mem_rdata_q[4] ;
 wire \mem_rdata_q[5] ;
 wire \mem_rdata_q[6] ;
 wire \mem_rdata_q[7] ;
 wire \mem_rdata_q[8] ;
 wire \mem_rdata_q[9] ;
 wire \mem_state[0] ;
 wire \mem_state[1] ;
 wire \mem_wordsize[0] ;
 wire \mem_wordsize[1] ;
 wire \mem_wordsize[2] ;
 wire pcpi_timeout;
 wire \pcpi_timeout_counter[0] ;
 wire \pcpi_timeout_counter[1] ;
 wire \pcpi_timeout_counter[2] ;
 wire \pcpi_timeout_counter[3] ;
 wire \reg_next_pc[0] ;
 wire \reg_next_pc[10] ;
 wire \reg_next_pc[11] ;
 wire \reg_next_pc[12] ;
 wire \reg_next_pc[13] ;
 wire \reg_next_pc[14] ;
 wire \reg_next_pc[15] ;
 wire \reg_next_pc[16] ;
 wire \reg_next_pc[17] ;
 wire \reg_next_pc[18] ;
 wire \reg_next_pc[19] ;
 wire \reg_next_pc[1] ;
 wire \reg_next_pc[20] ;
 wire \reg_next_pc[21] ;
 wire \reg_next_pc[22] ;
 wire \reg_next_pc[23] ;
 wire \reg_next_pc[24] ;
 wire \reg_next_pc[25] ;
 wire \reg_next_pc[26] ;
 wire \reg_next_pc[27] ;
 wire \reg_next_pc[28] ;
 wire \reg_next_pc[29] ;
 wire \reg_next_pc[2] ;
 wire \reg_next_pc[30] ;
 wire \reg_next_pc[31] ;
 wire \reg_next_pc[3] ;
 wire \reg_next_pc[4] ;
 wire \reg_next_pc[5] ;
 wire \reg_next_pc[6] ;
 wire \reg_next_pc[7] ;
 wire \reg_next_pc[8] ;
 wire \reg_next_pc[9] ;
 wire \reg_out[0] ;
 wire \reg_out[10] ;
 wire \reg_out[11] ;
 wire \reg_out[12] ;
 wire \reg_out[13] ;
 wire \reg_out[14] ;
 wire \reg_out[15] ;
 wire \reg_out[16] ;
 wire \reg_out[17] ;
 wire \reg_out[18] ;
 wire \reg_out[19] ;
 wire \reg_out[1] ;
 wire \reg_out[20] ;
 wire \reg_out[21] ;
 wire \reg_out[22] ;
 wire \reg_out[23] ;
 wire \reg_out[24] ;
 wire \reg_out[25] ;
 wire \reg_out[26] ;
 wire \reg_out[27] ;
 wire \reg_out[28] ;
 wire \reg_out[29] ;
 wire \reg_out[2] ;
 wire \reg_out[30] ;
 wire \reg_out[31] ;
 wire \reg_out[3] ;
 wire \reg_out[4] ;
 wire \reg_out[5] ;
 wire \reg_out[6] ;
 wire \reg_out[7] ;
 wire \reg_out[8] ;
 wire \reg_out[9] ;
 wire \reg_pc[10] ;
 wire \reg_pc[11] ;
 wire \reg_pc[12] ;
 wire \reg_pc[13] ;
 wire \reg_pc[14] ;
 wire \reg_pc[15] ;
 wire \reg_pc[16] ;
 wire \reg_pc[17] ;
 wire \reg_pc[18] ;
 wire \reg_pc[19] ;
 wire \reg_pc[1] ;
 wire \reg_pc[20] ;
 wire \reg_pc[21] ;
 wire \reg_pc[22] ;
 wire \reg_pc[23] ;
 wire \reg_pc[24] ;
 wire \reg_pc[25] ;
 wire \reg_pc[26] ;
 wire \reg_pc[27] ;
 wire \reg_pc[28] ;
 wire \reg_pc[29] ;
 wire \reg_pc[2] ;
 wire \reg_pc[30] ;
 wire \reg_pc[31] ;
 wire \reg_pc[3] ;
 wire \reg_pc[4] ;
 wire \reg_pc[5] ;
 wire \reg_pc[6] ;
 wire \reg_pc[7] ;
 wire \reg_pc[8] ;
 wire \reg_pc[9] ;
 wire \timer[0] ;
 wire \timer[10] ;
 wire \timer[11] ;
 wire \timer[12] ;
 wire \timer[13] ;
 wire \timer[14] ;
 wire \timer[15] ;
 wire \timer[16] ;
 wire \timer[17] ;
 wire \timer[18] ;
 wire \timer[19] ;
 wire \timer[1] ;
 wire \timer[20] ;
 wire \timer[21] ;
 wire \timer[22] ;
 wire \timer[23] ;
 wire \timer[24] ;
 wire \timer[25] ;
 wire \timer[26] ;
 wire \timer[27] ;
 wire \timer[28] ;
 wire \timer[29] ;
 wire \timer[2] ;
 wire \timer[30] ;
 wire \timer[31] ;
 wire \timer[3] ;
 wire \timer[4] ;
 wire \timer[5] ;
 wire \timer[6] ;
 wire \timer[7] ;
 wire \timer[8] ;
 wire \timer[9] ;
 wire net379;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net380;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net381;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire clknet_leaf_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;

 sky130_fd_sc_hd__clkbuf_2 _14652_ (.A(net66),
    .X(_08136_));
 sky130_fd_sc_hd__nand2_2 _14653_ (.A(net331),
    .B(_08136_),
    .Y(_08137_));
 sky130_fd_sc_hd__nand2_1 _14654_ (.A(net246),
    .B(net235),
    .Y(_08138_));
 sky130_fd_sc_hd__or4_1 _14655_ (.A(net260),
    .B(net257),
    .C(_08137_),
    .D(_08138_),
    .X(_08139_));
 sky130_fd_sc_hd__or3_1 _14656_ (.A(net256),
    .B(net259),
    .C(net240),
    .X(_08140_));
 sky130_fd_sc_hd__or4b_1 _14657_ (.A(net255),
    .B(net254),
    .C(net258),
    .D_N(net252),
    .X(_08141_));
 sky130_fd_sc_hd__or4bb_1 _14658_ (.A(net263),
    .B(net253),
    .C_N(net262),
    .D_N(net261),
    .X(_08142_));
 sky130_fd_sc_hd__or4_4 _14659_ (.A(_08139_),
    .B(_08140_),
    .C(_08141_),
    .D(_08142_),
    .X(_08143_));
 sky130_fd_sc_hd__o21ba_1 _14660_ (.A1(net239),
    .A2(net238),
    .B1_N(_08143_),
    .X(_08144_));
 sky130_fd_sc_hd__buf_1 _14661_ (.A(_08144_),
    .X(\genblk1.pcpi_mul.instr_any_mulh ));
 sky130_vsdinv _14662_ (.A(\cpu_state[1] ),
    .Y(_08145_));
 sky130_fd_sc_hd__clkbuf_2 _14663_ (.A(_08136_),
    .X(_08146_));
 sky130_fd_sc_hd__nand2_2 _14664_ (.A(_08145_),
    .B(_08146_),
    .Y(_08147_));
 sky130_fd_sc_hd__or2_4 _14665_ (.A(\cpu_state[5] ),
    .B(\cpu_state[6] ),
    .X(_08148_));
 sky130_fd_sc_hd__clkbuf_4 _14666_ (.A(_08148_),
    .X(_08149_));
 sky130_fd_sc_hd__or4_1 _14667_ (.A(instr_lb),
    .B(instr_lbu),
    .C(instr_lh),
    .D(instr_lhu),
    .X(_08150_));
 sky130_fd_sc_hd__clkbuf_2 _14668_ (.A(mem_do_rdata),
    .X(_08151_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14669_ (.A(\cpu_state[6] ),
    .X(_08152_));
 sky130_fd_sc_hd__clkbuf_2 _14670_ (.A(mem_do_prefetch),
    .X(_08153_));
 sky130_fd_sc_hd__nor2_1 _14671_ (.A(\mem_state[1] ),
    .B(\mem_state[0] ),
    .Y(_08154_));
 sky130_fd_sc_hd__nand2_2 _14672_ (.A(net65),
    .B(net198),
    .Y(_08155_));
 sky130_fd_sc_hd__and2_1 _14673_ (.A(\mem_state[1] ),
    .B(\mem_state[0] ),
    .X(_08156_));
 sky130_fd_sc_hd__a2bb2o_1 _14674_ (.A1_N(_08154_),
    .A2_N(_08155_),
    .B1(mem_do_rinst),
    .B2(_08156_),
    .X(_08157_));
 sky130_fd_sc_hd__o31a_1 _14675_ (.A1(mem_do_wdata),
    .A2(mem_do_rdata),
    .A3(mem_do_rinst),
    .B1(_08157_),
    .X(_08158_));
 sky130_fd_sc_hd__nand2_1 _14676_ (.A(_08136_),
    .B(_08158_),
    .Y(_08159_));
 sky130_fd_sc_hd__nand2_1 _14677_ (.A(_08153_),
    .B(_08159_),
    .Y(_08160_));
 sky130_fd_sc_hd__and4b_1 _14678_ (.A_N(_08151_),
    .B(_08136_),
    .C(_08152_),
    .D(_08160_),
    .X(_08161_));
 sky130_fd_sc_hd__or3b_1 _14679_ (.A(_08150_),
    .B(instr_lw),
    .C_N(_08161_),
    .X(_08162_));
 sky130_fd_sc_hd__clkbuf_2 _14680_ (.A(mem_do_wdata),
    .X(_08163_));
 sky130_fd_sc_hd__and4b_2 _14681_ (.A_N(_08163_),
    .B(_08136_),
    .C(\cpu_state[5] ),
    .D(_08160_),
    .X(_08164_));
 sky130_fd_sc_hd__or4b_1 _14682_ (.A(instr_sw),
    .B(instr_sh),
    .C(instr_sb),
    .D_N(_08164_),
    .X(_08165_));
 sky130_fd_sc_hd__o211a_1 _14683_ (.A1(_08147_),
    .A2(_08149_),
    .B1(_08162_),
    .C1(_08165_),
    .X(_08166_));
 sky130_fd_sc_hd__and2_1 _14684_ (.A(mem_do_prefetch),
    .B(_08159_),
    .X(_08167_));
 sky130_fd_sc_hd__o21a_1 _14685_ (.A1(_08151_),
    .A2(_08167_),
    .B1(\cpu_state[6] ),
    .X(_08168_));
 sky130_vsdinv _14686_ (.A(net66),
    .Y(_08169_));
 sky130_fd_sc_hd__clkbuf_2 _14687_ (.A(_08169_),
    .X(_08170_));
 sky130_fd_sc_hd__a311o_1 _14688_ (.A1(mem_do_wdata),
    .A2(\cpu_state[5] ),
    .A3(_08160_),
    .B1(_08168_),
    .C1(_08170_),
    .X(_08171_));
 sky130_fd_sc_hd__a21oi_4 _14689_ (.A1(\cpu_state[5] ),
    .A2(_08167_),
    .B1(_08171_),
    .Y(_08172_));
 sky130_fd_sc_hd__nand2_1 _14690_ (.A(_08166_),
    .B(_08172_),
    .Y(_08173_));
 sky130_fd_sc_hd__clkbuf_2 _14691_ (.A(_08161_),
    .X(_08174_));
 sky130_fd_sc_hd__nor2_2 _14692_ (.A(_08145_),
    .B(_08169_),
    .Y(_08175_));
 sky130_fd_sc_hd__clkbuf_4 _14693_ (.A(_08175_),
    .X(_08176_));
 sky130_fd_sc_hd__a221o_1 _14694_ (.A1(instr_sw),
    .A2(_08164_),
    .B1(_08174_),
    .B2(instr_lw),
    .C1(_08176_),
    .X(_08177_));
 sky130_fd_sc_hd__a21o_1 _14695_ (.A1(net459),
    .A2(_08173_),
    .B1(_08177_),
    .X(_00047_));
 sky130_fd_sc_hd__clkbuf_4 _14696_ (.A(\cpu_state[2] ),
    .X(_08178_));
 sky130_fd_sc_hd__clkbuf_2 _14697_ (.A(_08178_),
    .X(_08179_));
 sky130_fd_sc_hd__clkbuf_2 _14698_ (.A(_08179_),
    .X(_08180_));
 sky130_fd_sc_hd__clkbuf_2 _14699_ (.A(_08180_),
    .X(_08181_));
 sky130_fd_sc_hd__buf_2 _14700_ (.A(_08170_),
    .X(_08182_));
 sky130_fd_sc_hd__buf_2 _14701_ (.A(_08182_),
    .X(_08183_));
 sky130_fd_sc_hd__buf_2 _14702_ (.A(\reg_pc[1] ),
    .X(_08184_));
 sky130_fd_sc_hd__o21a_1 _14703_ (.A1(\reg_next_pc[0] ),
    .A2(_08184_),
    .B1(mem_do_rinst),
    .X(_08185_));
 sky130_fd_sc_hd__clkbuf_2 _14704_ (.A(irq_active),
    .X(_08186_));
 sky130_fd_sc_hd__nor2_1 _14705_ (.A(\irq_mask[2] ),
    .B(_08186_),
    .Y(_08187_));
 sky130_fd_sc_hd__and3_1 _14706_ (.A(_08136_),
    .B(_08185_),
    .C(_08187_),
    .X(_08188_));
 sky130_vsdinv _14707_ (.A(_08185_),
    .Y(_08189_));
 sky130_fd_sc_hd__nor2_1 _14708_ (.A(_08170_),
    .B(_08189_),
    .Y(_08190_));
 sky130_fd_sc_hd__clkbuf_2 _14709_ (.A(net267),
    .X(_08191_));
 sky130_fd_sc_hd__nand2_1 _14710_ (.A(\mem_wordsize[2] ),
    .B(_08191_),
    .Y(_08192_));
 sky130_fd_sc_hd__buf_2 _14711_ (.A(net278),
    .X(_08193_));
 sky130_fd_sc_hd__o21ai_2 _14712_ (.A1(net267),
    .A2(_08193_),
    .B1(\mem_wordsize[0] ),
    .Y(_08194_));
 sky130_fd_sc_hd__nand2_1 _14713_ (.A(_08192_),
    .B(_08194_),
    .Y(_08195_));
 sky130_fd_sc_hd__nor2_1 _14714_ (.A(_08190_),
    .B(_08195_),
    .Y(_08196_));
 sky130_fd_sc_hd__nor2_1 _14715_ (.A(mem_do_wdata),
    .B(mem_do_rdata),
    .Y(_08197_));
 sky130_fd_sc_hd__nor2_1 _14716_ (.A(_08170_),
    .B(_08197_),
    .Y(_08198_));
 sky130_fd_sc_hd__and3b_1 _14717_ (.A_N(_08192_),
    .B(_08187_),
    .C(_08198_),
    .X(_08199_));
 sky130_fd_sc_hd__nor2_1 _14718_ (.A(_08190_),
    .B(_08198_),
    .Y(_08200_));
 sky130_fd_sc_hd__and4b_1 _14719_ (.A_N(_08194_),
    .B(_08187_),
    .C(_08198_),
    .D(_08192_),
    .X(_08201_));
 sky130_fd_sc_hd__and2b_1 _14720_ (.A_N(_08190_),
    .B(_08201_),
    .X(_08202_));
 sky130_fd_sc_hd__a211o_1 _14721_ (.A1(_08189_),
    .A2(_08199_),
    .B1(_08200_),
    .C1(_08202_),
    .X(_08203_));
 sky130_fd_sc_hd__or3_2 _14722_ (.A(_08188_),
    .B(_08196_),
    .C(_08203_),
    .X(_08204_));
 sky130_vsdinv _14723_ (.A(_08204_),
    .Y(_08205_));
 sky130_fd_sc_hd__nor2_2 _14724_ (.A(_08183_),
    .B(_08205_),
    .Y(_08206_));
 sky130_fd_sc_hd__clkbuf_4 _14725_ (.A(instr_waitirq),
    .X(_08207_));
 sky130_fd_sc_hd__or3_1 _14726_ (.A(instr_sw),
    .B(instr_sh),
    .C(instr_sb),
    .X(_08208_));
 sky130_fd_sc_hd__or4_1 _14727_ (.A(_08207_),
    .B(instr_slli),
    .C(instr_jalr),
    .D(_08208_),
    .X(_08209_));
 sky130_fd_sc_hd__or4_1 _14728_ (.A(instr_bltu),
    .B(instr_blt),
    .C(instr_bne),
    .D(instr_beq),
    .X(_08210_));
 sky130_fd_sc_hd__or4_1 _14729_ (.A(instr_andi),
    .B(instr_ori),
    .C(instr_xori),
    .D(_08210_),
    .X(_08211_));
 sky130_fd_sc_hd__or4_1 _14730_ (.A(instr_and),
    .B(instr_or),
    .C(instr_bgeu),
    .D(instr_bge),
    .X(_08212_));
 sky130_fd_sc_hd__or4_1 _14731_ (.A(instr_xor),
    .B(instr_sll),
    .C(instr_sub),
    .D(instr_add),
    .X(_08213_));
 sky130_fd_sc_hd__or4_1 _14732_ (.A(instr_lw),
    .B(_08150_),
    .C(_08212_),
    .D(_08213_),
    .X(_08214_));
 sky130_fd_sc_hd__or4_1 _14733_ (.A(instr_addi),
    .B(_08209_),
    .C(_08211_),
    .D(_08214_),
    .X(_08215_));
 sky130_fd_sc_hd__or2_2 _14734_ (.A(instr_auipc),
    .B(instr_lui),
    .X(_08216_));
 sky130_fd_sc_hd__or2_1 _14735_ (.A(instr_jal),
    .B(_08216_),
    .X(_08217_));
 sky130_fd_sc_hd__clkbuf_2 _14736_ (.A(_08217_),
    .X(_00037_));
 sky130_fd_sc_hd__or4_2 _14737_ (.A(instr_sra),
    .B(instr_srl),
    .C(instr_srli),
    .D(instr_srai),
    .X(_08218_));
 sky130_fd_sc_hd__or4_1 _14738_ (.A(instr_sltu),
    .B(instr_slt),
    .C(instr_sltiu),
    .D(instr_slti),
    .X(_08219_));
 sky130_fd_sc_hd__or3_1 _14739_ (.A(_00037_),
    .B(_08218_),
    .C(_08219_),
    .X(_08220_));
 sky130_fd_sc_hd__nor3_1 _14740_ (.A(instr_retirq),
    .B(instr_getq),
    .C(instr_setq),
    .Y(_08221_));
 sky130_fd_sc_hd__or3b_1 _14741_ (.A(instr_timer),
    .B(instr_maskirq),
    .C_N(_08221_),
    .X(_08222_));
 sky130_fd_sc_hd__nor3_1 _14742_ (.A(instr_rdinstr),
    .B(instr_rdinstrh),
    .C(instr_rdcycleh),
    .Y(_08223_));
 sky130_fd_sc_hd__or3b_4 _14743_ (.A(instr_rdcycle),
    .B(_08222_),
    .C_N(_08223_),
    .X(_08224_));
 sky130_fd_sc_hd__nor3_1 _14744_ (.A(_08215_),
    .B(_08220_),
    .C(_08224_),
    .Y(_08225_));
 sky130_fd_sc_hd__or2b_1 _14745_ (.A(net369),
    .B_N(is_lb_lh_lw_lbu_lhu),
    .X(_08226_));
 sky130_vsdinv _14746_ (.A(_08226_),
    .Y(_08227_));
 sky130_vsdinv _14747_ (.A(_08158_),
    .Y(_08228_));
 sky130_fd_sc_hd__o21a_1 _14748_ (.A1(_08153_),
    .A2(_08228_),
    .B1(_08206_),
    .X(_08229_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14749_ (.A(_08152_),
    .X(_08230_));
 sky130_fd_sc_hd__clkbuf_2 _14750_ (.A(_08230_),
    .X(_08231_));
 sky130_fd_sc_hd__a32o_1 _14751_ (.A1(_08181_),
    .A2(_08206_),
    .A3(_08227_),
    .B1(_08229_),
    .B2(_08231_),
    .X(_00046_));
 sky130_fd_sc_hd__clkbuf_2 _14752_ (.A(\cpu_state[1] ),
    .X(_08232_));
 sky130_vsdinv _14753_ (.A(decoder_trigger),
    .Y(_08233_));
 sky130_fd_sc_hd__and2b_1 _14754_ (.A_N(\irq_mask[18] ),
    .B(\irq_pending[18] ),
    .X(_08234_));
 sky130_fd_sc_hd__and2b_2 _14755_ (.A_N(\irq_mask[11] ),
    .B(\irq_pending[11] ),
    .X(_08235_));
 sky130_fd_sc_hd__and2b_2 _14756_ (.A_N(\irq_mask[3] ),
    .B(\irq_pending[3] ),
    .X(_08236_));
 sky130_fd_sc_hd__and2b_2 _14757_ (.A_N(\irq_mask[8] ),
    .B(\irq_pending[8] ),
    .X(_08237_));
 sky130_fd_sc_hd__or4_1 _14758_ (.A(_08234_),
    .B(_08235_),
    .C(_08236_),
    .D(_08237_),
    .X(_08238_));
 sky130_fd_sc_hd__and2b_2 _14759_ (.A_N(\irq_mask[25] ),
    .B(\irq_pending[25] ),
    .X(_08239_));
 sky130_fd_sc_hd__and2b_2 _14760_ (.A_N(\irq_mask[0] ),
    .B(\irq_pending[0] ),
    .X(_08240_));
 sky130_fd_sc_hd__and2b_2 _14761_ (.A_N(\irq_mask[26] ),
    .B(\irq_pending[26] ),
    .X(_08241_));
 sky130_fd_sc_hd__and2b_2 _14762_ (.A_N(\irq_mask[29] ),
    .B(\irq_pending[29] ),
    .X(_08242_));
 sky130_fd_sc_hd__or4_1 _14763_ (.A(_08239_),
    .B(_08240_),
    .C(_08241_),
    .D(_08242_),
    .X(_08243_));
 sky130_fd_sc_hd__and2b_2 _14764_ (.A_N(\irq_mask[20] ),
    .B(\irq_pending[20] ),
    .X(_08244_));
 sky130_fd_sc_hd__and2b_2 _14765_ (.A_N(\irq_mask[22] ),
    .B(\irq_pending[22] ),
    .X(_08245_));
 sky130_fd_sc_hd__and2b_2 _14766_ (.A_N(\irq_mask[21] ),
    .B(\irq_pending[21] ),
    .X(_08246_));
 sky130_fd_sc_hd__and2b_2 _14767_ (.A_N(\irq_mask[10] ),
    .B(\irq_pending[10] ),
    .X(_08247_));
 sky130_fd_sc_hd__or4_1 _14768_ (.A(_08244_),
    .B(_08245_),
    .C(_08246_),
    .D(_08247_),
    .X(_08248_));
 sky130_fd_sc_hd__and2b_2 _14769_ (.A_N(\irq_mask[23] ),
    .B(\irq_pending[23] ),
    .X(_08249_));
 sky130_fd_sc_hd__and2b_2 _14770_ (.A_N(\irq_mask[15] ),
    .B(\irq_pending[15] ),
    .X(_08250_));
 sky130_fd_sc_hd__and2b_2 _14771_ (.A_N(\irq_mask[12] ),
    .B(\irq_pending[12] ),
    .X(_08251_));
 sky130_fd_sc_hd__and2b_2 _14772_ (.A_N(\irq_mask[9] ),
    .B(\irq_pending[9] ),
    .X(_08252_));
 sky130_fd_sc_hd__or4_1 _14773_ (.A(_08249_),
    .B(_08250_),
    .C(_08251_),
    .D(_08252_),
    .X(_08253_));
 sky130_fd_sc_hd__or4_1 _14774_ (.A(_08238_),
    .B(_08243_),
    .C(_08248_),
    .D(_08253_),
    .X(_08254_));
 sky130_fd_sc_hd__and2b_2 _14775_ (.A_N(\irq_mask[19] ),
    .B(\irq_pending[19] ),
    .X(_08255_));
 sky130_fd_sc_hd__and2b_2 _14776_ (.A_N(\irq_mask[28] ),
    .B(\irq_pending[28] ),
    .X(_08256_));
 sky130_fd_sc_hd__and2b_2 _14777_ (.A_N(\irq_mask[16] ),
    .B(\irq_pending[16] ),
    .X(_08257_));
 sky130_fd_sc_hd__and2b_2 _14778_ (.A_N(\irq_mask[31] ),
    .B(\irq_pending[31] ),
    .X(_08258_));
 sky130_fd_sc_hd__or4_1 _14779_ (.A(_08255_),
    .B(_08256_),
    .C(_08257_),
    .D(_08258_),
    .X(_08259_));
 sky130_fd_sc_hd__and2b_2 _14780_ (.A_N(\irq_mask[13] ),
    .B(\irq_pending[13] ),
    .X(_08260_));
 sky130_fd_sc_hd__and2b_2 _14781_ (.A_N(\irq_mask[27] ),
    .B(\irq_pending[27] ),
    .X(_08261_));
 sky130_fd_sc_hd__and2b_2 _14782_ (.A_N(\irq_mask[24] ),
    .B(\irq_pending[24] ),
    .X(_08262_));
 sky130_fd_sc_hd__and2b_2 _14783_ (.A_N(\irq_mask[1] ),
    .B(\irq_pending[1] ),
    .X(_08263_));
 sky130_fd_sc_hd__or4_1 _14784_ (.A(_08260_),
    .B(_08261_),
    .C(_08262_),
    .D(_08263_),
    .X(_08264_));
 sky130_fd_sc_hd__and2b_2 _14785_ (.A_N(\irq_mask[5] ),
    .B(\irq_pending[5] ),
    .X(_08265_));
 sky130_fd_sc_hd__and2b_2 _14786_ (.A_N(\irq_mask[6] ),
    .B(\irq_pending[6] ),
    .X(_08266_));
 sky130_fd_sc_hd__and2b_2 _14787_ (.A_N(\irq_mask[4] ),
    .B(\irq_pending[4] ),
    .X(_08267_));
 sky130_fd_sc_hd__and2b_2 _14788_ (.A_N(\irq_mask[2] ),
    .B(\irq_pending[2] ),
    .X(_08268_));
 sky130_fd_sc_hd__or4_1 _14789_ (.A(_08265_),
    .B(_08266_),
    .C(_08267_),
    .D(_08268_),
    .X(_08269_));
 sky130_fd_sc_hd__and2b_2 _14790_ (.A_N(\irq_mask[30] ),
    .B(\irq_pending[30] ),
    .X(_08270_));
 sky130_fd_sc_hd__and2b_2 _14791_ (.A_N(\irq_mask[14] ),
    .B(\irq_pending[14] ),
    .X(_08271_));
 sky130_fd_sc_hd__and2b_2 _14792_ (.A_N(\irq_mask[17] ),
    .B(\irq_pending[17] ),
    .X(_08272_));
 sky130_fd_sc_hd__and2b_2 _14793_ (.A_N(\irq_mask[7] ),
    .B(\irq_pending[7] ),
    .X(_08273_));
 sky130_fd_sc_hd__or4_1 _14794_ (.A(_08270_),
    .B(_08271_),
    .C(_08272_),
    .D(_08273_),
    .X(_08274_));
 sky130_fd_sc_hd__or4_1 _14795_ (.A(_08259_),
    .B(_08264_),
    .C(_08269_),
    .D(_08274_),
    .X(_08275_));
 sky130_fd_sc_hd__nor2_1 _14796_ (.A(irq_active),
    .B(irq_delay),
    .Y(_08276_));
 sky130_fd_sc_hd__o211a_1 _14797_ (.A1(_08254_),
    .A2(_08275_),
    .B1(_08276_),
    .C1(decoder_trigger),
    .X(_08277_));
 sky130_fd_sc_hd__or2_4 _14798_ (.A(\irq_state[1] ),
    .B(\irq_state[0] ),
    .X(_08278_));
 sky130_fd_sc_hd__or4_4 _14799_ (.A(instr_waitirq),
    .B(_08233_),
    .C(_08277_),
    .D(_08278_),
    .X(_08279_));
 sky130_fd_sc_hd__clkbuf_2 _14800_ (.A(_08279_),
    .X(_08280_));
 sky130_fd_sc_hd__clkbuf_2 _14801_ (.A(\irq_mask[1] ),
    .X(_08281_));
 sky130_fd_sc_hd__nor2_1 _14802_ (.A(instr_ecall_ebreak),
    .B(pcpi_timeout),
    .Y(_08282_));
 sky130_fd_sc_hd__nor3_1 _14803_ (.A(_08281_),
    .B(_08186_),
    .C(_08282_),
    .Y(_08283_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14804_ (.A(\cpu_state[3] ),
    .X(_08284_));
 sky130_fd_sc_hd__buf_2 _14805_ (.A(_08284_),
    .X(_08285_));
 sky130_fd_sc_hd__buf_2 _14806_ (.A(_08285_),
    .X(_08286_));
 sky130_fd_sc_hd__clkbuf_2 _14807_ (.A(_08286_),
    .X(_08287_));
 sky130_fd_sc_hd__clkbuf_2 _14808_ (.A(_08287_),
    .X(_08288_));
 sky130_fd_sc_hd__o211a_1 _14809_ (.A1(\genblk1.pcpi_mul.active[1] ),
    .A2(_08283_),
    .B1(net369),
    .C1(_08288_),
    .X(_08289_));
 sky130_fd_sc_hd__nor2_1 _14810_ (.A(\cpu_state[5] ),
    .B(\cpu_state[6] ),
    .Y(_08290_));
 sky130_fd_sc_hd__buf_2 _14811_ (.A(_08290_),
    .X(_08291_));
 sky130_fd_sc_hd__or3_1 _14812_ (.A(_08153_),
    .B(_08159_),
    .C(_08291_),
    .X(_08292_));
 sky130_fd_sc_hd__inv_2 _14813_ (.A(_08292_),
    .Y(_01169_));
 sky130_fd_sc_hd__clkbuf_2 _14814_ (.A(_08179_),
    .X(_08293_));
 sky130_fd_sc_hd__buf_2 _14815_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_08294_));
 sky130_vsdinv _14816_ (.A(\cpu_state[4] ),
    .Y(_08295_));
 sky130_fd_sc_hd__or2_1 _14817_ (.A(_08295_),
    .B(alu_wait),
    .X(_08296_));
 sky130_fd_sc_hd__nor2_1 _14818_ (.A(_08294_),
    .B(_08296_),
    .Y(_08297_));
 sky130_fd_sc_hd__a21o_1 _14819_ (.A1(_08293_),
    .A2(_08224_),
    .B1(_08297_),
    .X(_08298_));
 sky130_fd_sc_hd__a2111o_1 _14820_ (.A1(_08232_),
    .A2(_08280_),
    .B1(_08289_),
    .C1(_01169_),
    .D1(_08298_),
    .X(_08299_));
 sky130_fd_sc_hd__or2_1 _14821_ (.A(_08182_),
    .B(_08197_),
    .X(_08300_));
 sky130_fd_sc_hd__nor4_1 _14822_ (.A(_08202_),
    .B(_08188_),
    .C(_08200_),
    .D(_08199_),
    .Y(_08301_));
 sky130_fd_sc_hd__o21ai_1 _14823_ (.A1(_08300_),
    .A2(_08195_),
    .B1(net368),
    .Y(_08302_));
 sky130_vsdinv _14824_ (.A(instr_jal),
    .Y(_08303_));
 sky130_fd_sc_hd__nor2_2 _14825_ (.A(_08303_),
    .B(_08233_),
    .Y(_08304_));
 sky130_fd_sc_hd__or2_1 _14826_ (.A(decoder_trigger),
    .B(do_waitirq),
    .X(_08305_));
 sky130_fd_sc_hd__and2_2 _14827_ (.A(_08207_),
    .B(_08305_),
    .X(_08306_));
 sky130_fd_sc_hd__or2_2 _14828_ (.A(_08277_),
    .B(_08278_),
    .X(_08307_));
 sky130_fd_sc_hd__nor2_2 _14829_ (.A(_08306_),
    .B(_08307_),
    .Y(_08308_));
 sky130_fd_sc_hd__clkbuf_4 _14830_ (.A(_08308_),
    .X(_08309_));
 sky130_fd_sc_hd__a21boi_1 _14831_ (.A1(_08185_),
    .A2(net368),
    .B1_N(_08309_),
    .Y(_08310_));
 sky130_fd_sc_hd__clkbuf_2 _14832_ (.A(\cpu_state[4] ),
    .X(_08311_));
 sky130_fd_sc_hd__clkbuf_2 _14833_ (.A(_08311_),
    .X(_08312_));
 sky130_vsdinv _14834_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .Y(_08313_));
 sky130_fd_sc_hd__nor2_1 _14835_ (.A(_08313_),
    .B(alu_wait),
    .Y(_08314_));
 sky130_fd_sc_hd__and2_1 _14836_ (.A(_08312_),
    .B(_08314_),
    .X(_08315_));
 sky130_fd_sc_hd__a31o_1 _14837_ (.A1(_08158_),
    .A2(_08204_),
    .A3(_08315_),
    .B1(_08183_),
    .X(_08316_));
 sky130_fd_sc_hd__a41o_1 _14838_ (.A1(_08232_),
    .A2(_08302_),
    .A3(_08304_),
    .A4(_08310_),
    .B1(_08316_),
    .X(_08317_));
 sky130_fd_sc_hd__a21o_1 _14839_ (.A1(_08204_),
    .A2(_08299_),
    .B1(_08317_),
    .X(_00041_));
 sky130_fd_sc_hd__nand2_1 _14840_ (.A(_08286_),
    .B(net369),
    .Y(_08318_));
 sky130_fd_sc_hd__or2_1 _14841_ (.A(\genblk1.pcpi_mul.active[1] ),
    .B(_08318_),
    .X(_08319_));
 sky130_vsdinv _14842_ (.A(_08319_),
    .Y(_08320_));
 sky130_fd_sc_hd__buf_2 _14843_ (.A(_08146_),
    .X(_08321_));
 sky130_fd_sc_hd__clkbuf_4 _14844_ (.A(_08321_),
    .X(_08322_));
 sky130_fd_sc_hd__o221a_1 _14845_ (.A1(_08281_),
    .A2(_08186_),
    .B1(instr_ecall_ebreak),
    .B2(pcpi_timeout),
    .C1(_08322_),
    .X(_08323_));
 sky130_fd_sc_hd__buf_2 _14846_ (.A(\mem_wordsize[2] ),
    .X(_08324_));
 sky130_fd_sc_hd__buf_2 _14847_ (.A(_08191_),
    .X(_08325_));
 sky130_fd_sc_hd__buf_2 _14848_ (.A(_08325_),
    .X(_08326_));
 sky130_fd_sc_hd__a31o_1 _14849_ (.A1(_08324_),
    .A2(_08326_),
    .A3(_08187_),
    .B1(_08197_),
    .X(_08327_));
 sky130_fd_sc_hd__clkbuf_2 _14850_ (.A(_08146_),
    .X(_08328_));
 sky130_fd_sc_hd__a2bb2o_1 _14851_ (.A1_N(_08300_),
    .A2_N(_08195_),
    .B1(_08327_),
    .B2(_08328_),
    .X(_08329_));
 sky130_fd_sc_hd__o31a_1 _14852_ (.A1(_08190_),
    .A2(_08201_),
    .A3(_08329_),
    .B1(\cpu_state[0] ),
    .X(_08330_));
 sky130_fd_sc_hd__a211o_1 _14853_ (.A1(_08320_),
    .A2(_08323_),
    .B1(_08330_),
    .C1(_08205_),
    .X(_00040_));
 sky130_fd_sc_hd__clkbuf_2 _14854_ (.A(_08308_),
    .X(_08331_));
 sky130_fd_sc_hd__clkbuf_4 _14855_ (.A(_08331_),
    .X(_08332_));
 sky130_fd_sc_hd__nand2_1 _14856_ (.A(_08207_),
    .B(_08305_),
    .Y(_08333_));
 sky130_fd_sc_hd__clkbuf_4 _14857_ (.A(_08333_),
    .X(_08334_));
 sky130_fd_sc_hd__a21bo_1 _14858_ (.A1(_08187_),
    .A2(_08334_),
    .B1_N(_08190_),
    .X(_08335_));
 sky130_fd_sc_hd__clkbuf_2 _14859_ (.A(instr_jal),
    .X(_08336_));
 sky130_fd_sc_hd__nor2_1 _14860_ (.A(_08336_),
    .B(_08233_),
    .Y(_08337_));
 sky130_fd_sc_hd__buf_2 _14861_ (.A(_08337_),
    .X(_08338_));
 sky130_fd_sc_hd__and3_1 _14862_ (.A(_08176_),
    .B(_08335_),
    .C(_08338_),
    .X(_08339_));
 sky130_fd_sc_hd__and3_1 _14863_ (.A(_08332_),
    .B(_08302_),
    .C(_08339_),
    .X(_08340_));
 sky130_fd_sc_hd__clkbuf_1 _14864_ (.A(_08340_),
    .X(_00042_));
 sky130_fd_sc_hd__and2_1 _14865_ (.A(net270),
    .B(net302),
    .X(_08341_));
 sky130_fd_sc_hd__clkbuf_2 _14866_ (.A(net270),
    .X(_08342_));
 sky130_fd_sc_hd__clkbuf_4 _14867_ (.A(net302),
    .X(_08343_));
 sky130_fd_sc_hd__nor2_1 _14868_ (.A(_08342_),
    .B(_08343_),
    .Y(_08344_));
 sky130_fd_sc_hd__nor2_2 _14869_ (.A(_08341_),
    .B(_08344_),
    .Y(_08345_));
 sky130_fd_sc_hd__clkbuf_2 _14870_ (.A(net271),
    .X(_08346_));
 sky130_fd_sc_hd__clkbuf_4 _14871_ (.A(net303),
    .X(_08347_));
 sky130_fd_sc_hd__nor2_1 _14872_ (.A(_08346_),
    .B(_08347_),
    .Y(_08348_));
 sky130_fd_sc_hd__and2_1 _14873_ (.A(_08346_),
    .B(net303),
    .X(_08349_));
 sky130_fd_sc_hd__nor2_2 _14874_ (.A(_08348_),
    .B(_08349_),
    .Y(_08350_));
 sky130_fd_sc_hd__clkbuf_2 _14875_ (.A(net276),
    .X(_08351_));
 sky130_fd_sc_hd__and2_1 _14876_ (.A(_08351_),
    .B(net308),
    .X(_08352_));
 sky130_fd_sc_hd__nor2_1 _14877_ (.A(_08351_),
    .B(net308),
    .Y(_08353_));
 sky130_fd_sc_hd__nor2_1 _14878_ (.A(_08352_),
    .B(_08353_),
    .Y(_08354_));
 sky130_fd_sc_hd__clkbuf_2 _14879_ (.A(net279),
    .X(_08355_));
 sky130_fd_sc_hd__and2_1 _14880_ (.A(_08355_),
    .B(net311),
    .X(_08356_));
 sky130_fd_sc_hd__nor2_1 _14881_ (.A(_08355_),
    .B(net311),
    .Y(_08357_));
 sky130_fd_sc_hd__nor2_1 _14882_ (.A(_08356_),
    .B(_08357_),
    .Y(_08358_));
 sky130_fd_sc_hd__clkbuf_2 _14883_ (.A(net281),
    .X(_08359_));
 sky130_fd_sc_hd__and2_1 _14884_ (.A(_08359_),
    .B(net313),
    .X(_08360_));
 sky130_fd_sc_hd__nor2_1 _14885_ (.A(_08359_),
    .B(net313),
    .Y(_08361_));
 sky130_fd_sc_hd__nor2_1 _14886_ (.A(_08360_),
    .B(_08361_),
    .Y(_08362_));
 sky130_fd_sc_hd__clkbuf_2 _14887_ (.A(net280),
    .X(_08363_));
 sky130_fd_sc_hd__clkbuf_2 _14888_ (.A(net312),
    .X(_08364_));
 sky130_fd_sc_hd__nor2_1 _14889_ (.A(_08363_),
    .B(_08364_),
    .Y(_08365_));
 sky130_fd_sc_hd__nand2_1 _14890_ (.A(net280),
    .B(net312),
    .Y(_08366_));
 sky130_fd_sc_hd__nor2b_2 _14891_ (.A(_08365_),
    .B_N(_08366_),
    .Y(_08367_));
 sky130_fd_sc_hd__nor2_1 _14892_ (.A(net282),
    .B(net314),
    .Y(_08368_));
 sky130_fd_sc_hd__buf_2 _14893_ (.A(net314),
    .X(_08369_));
 sky130_fd_sc_hd__nand2_1 _14894_ (.A(net282),
    .B(_08369_),
    .Y(_08370_));
 sky130_fd_sc_hd__and2b_1 _14895_ (.A_N(_08368_),
    .B(_08370_),
    .X(_08371_));
 sky130_fd_sc_hd__or4_1 _14896_ (.A(_08358_),
    .B(_08362_),
    .C(_08367_),
    .D(_08371_),
    .X(_08372_));
 sky130_fd_sc_hd__nor2_1 _14897_ (.A(net277),
    .B(net309),
    .Y(_08373_));
 sky130_fd_sc_hd__clkbuf_2 _14898_ (.A(net277),
    .X(_08374_));
 sky130_fd_sc_hd__clkbuf_4 _14899_ (.A(net309),
    .X(_08375_));
 sky130_fd_sc_hd__nand2_1 _14900_ (.A(_08374_),
    .B(_08375_),
    .Y(_08376_));
 sky130_fd_sc_hd__nor2b_2 _14901_ (.A(_08373_),
    .B_N(_08376_),
    .Y(_08377_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14902_ (.A(net274),
    .X(_08378_));
 sky130_fd_sc_hd__and2_1 _14903_ (.A(_08378_),
    .B(net306),
    .X(_08379_));
 sky130_fd_sc_hd__nor2_1 _14904_ (.A(_08378_),
    .B(net306),
    .Y(_08380_));
 sky130_fd_sc_hd__nor2_1 _14905_ (.A(_08379_),
    .B(_08380_),
    .Y(_08381_));
 sky130_fd_sc_hd__buf_1 _14906_ (.A(net275),
    .X(_08382_));
 sky130_fd_sc_hd__clkbuf_4 _14907_ (.A(net307),
    .X(_08383_));
 sky130_fd_sc_hd__or2_1 _14908_ (.A(_08382_),
    .B(_08383_),
    .X(_08384_));
 sky130_fd_sc_hd__nand2_1 _14909_ (.A(net275),
    .B(net307),
    .Y(_08385_));
 sky130_fd_sc_hd__and2_1 _14910_ (.A(_08384_),
    .B(_08385_),
    .X(_08386_));
 sky130_fd_sc_hd__or2_1 _14911_ (.A(_08381_),
    .B(_08386_),
    .X(_08387_));
 sky130_fd_sc_hd__or4_1 _14912_ (.A(_08354_),
    .B(_08372_),
    .C(_08377_),
    .D(_08387_),
    .X(_08388_));
 sky130_fd_sc_hd__nor2_1 _14913_ (.A(net298),
    .B(net330),
    .Y(_08389_));
 sky130_fd_sc_hd__nand2_1 _14914_ (.A(net298),
    .B(net330),
    .Y(_08390_));
 sky130_fd_sc_hd__and2b_1 _14915_ (.A_N(_08389_),
    .B(_08390_),
    .X(_08391_));
 sky130_fd_sc_hd__or2_1 _14916_ (.A(net291),
    .B(net323),
    .X(_08392_));
 sky130_fd_sc_hd__buf_2 _14917_ (.A(net291),
    .X(_08393_));
 sky130_fd_sc_hd__nand2_1 _14918_ (.A(_08393_),
    .B(net323),
    .Y(_08394_));
 sky130_fd_sc_hd__and2_1 _14919_ (.A(_08392_),
    .B(_08394_),
    .X(_08395_));
 sky130_fd_sc_hd__or2_1 _14920_ (.A(net288),
    .B(net320),
    .X(_08396_));
 sky130_fd_sc_hd__clkbuf_2 _14921_ (.A(net288),
    .X(_08397_));
 sky130_fd_sc_hd__clkbuf_4 _14922_ (.A(net320),
    .X(_08398_));
 sky130_fd_sc_hd__nand2_1 _14923_ (.A(_08397_),
    .B(_08398_),
    .Y(_08399_));
 sky130_fd_sc_hd__and2_1 _14924_ (.A(_08396_),
    .B(_08399_),
    .X(_08400_));
 sky130_fd_sc_hd__clkbuf_2 _14925_ (.A(net268),
    .X(_08401_));
 sky130_fd_sc_hd__nand2_1 _14926_ (.A(_08401_),
    .B(net300),
    .Y(_08402_));
 sky130_fd_sc_hd__or2_1 _14927_ (.A(net268),
    .B(net300),
    .X(_08403_));
 sky130_fd_sc_hd__and2_1 _14928_ (.A(_08402_),
    .B(_08403_),
    .X(_08404_));
 sky130_fd_sc_hd__or4_1 _14929_ (.A(_08391_),
    .B(_08395_),
    .C(_08400_),
    .D(_08404_),
    .X(_08405_));
 sky130_fd_sc_hd__or4_1 _14930_ (.A(_08345_),
    .B(_08350_),
    .C(_08388_),
    .D(_08405_),
    .X(_08406_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14931_ (.A(net295),
    .X(_08407_));
 sky130_fd_sc_hd__or2_1 _14932_ (.A(net189),
    .B(_08407_),
    .X(_08408_));
 sky130_fd_sc_hd__nand2_1 _14933_ (.A(net189),
    .B(_08407_),
    .Y(_08409_));
 sky130_fd_sc_hd__and2_1 _14934_ (.A(_08408_),
    .B(_08409_),
    .X(_08410_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14935_ (.A(net269),
    .X(_08411_));
 sky130_fd_sc_hd__clkbuf_4 _14936_ (.A(_08411_),
    .X(_08412_));
 sky130_fd_sc_hd__clkbuf_4 _14937_ (.A(net301),
    .X(_08413_));
 sky130_fd_sc_hd__and2_1 _14938_ (.A(_08412_),
    .B(_08413_),
    .X(_08414_));
 sky130_fd_sc_hd__nor2_1 _14939_ (.A(net269),
    .B(net301),
    .Y(_08415_));
 sky130_fd_sc_hd__nor2_1 _14940_ (.A(_08414_),
    .B(_08415_),
    .Y(_08416_));
 sky130_fd_sc_hd__clkbuf_2 _14941_ (.A(net272),
    .X(_08417_));
 sky130_fd_sc_hd__and2_1 _14942_ (.A(_08417_),
    .B(net304),
    .X(_08418_));
 sky130_fd_sc_hd__clkbuf_4 _14943_ (.A(net304),
    .X(_08419_));
 sky130_fd_sc_hd__nor2_1 _14944_ (.A(_08417_),
    .B(_08419_),
    .Y(_08420_));
 sky130_fd_sc_hd__nor2_2 _14945_ (.A(_08418_),
    .B(_08420_),
    .Y(_08421_));
 sky130_fd_sc_hd__or3_1 _14946_ (.A(_08410_),
    .B(_08416_),
    .C(_08421_),
    .X(_08422_));
 sky130_fd_sc_hd__clkbuf_2 _14947_ (.A(net283),
    .X(_08423_));
 sky130_fd_sc_hd__and2_1 _14948_ (.A(_08423_),
    .B(net315),
    .X(_08424_));
 sky130_fd_sc_hd__nor2_1 _14949_ (.A(_08423_),
    .B(net315),
    .Y(_08425_));
 sky130_fd_sc_hd__nor2_2 _14950_ (.A(_08424_),
    .B(_08425_),
    .Y(_08426_));
 sky130_fd_sc_hd__clkbuf_4 _14951_ (.A(net316),
    .X(_08427_));
 sky130_fd_sc_hd__nor2_1 _14952_ (.A(net284),
    .B(_08427_),
    .Y(_08428_));
 sky130_fd_sc_hd__and2_1 _14953_ (.A(net284),
    .B(net316),
    .X(_08429_));
 sky130_fd_sc_hd__nor2_2 _14954_ (.A(_08428_),
    .B(_08429_),
    .Y(_08430_));
 sky130_fd_sc_hd__and2_1 _14955_ (.A(net285),
    .B(net317),
    .X(_08431_));
 sky130_fd_sc_hd__nor2_1 _14956_ (.A(net285),
    .B(net317),
    .Y(_08432_));
 sky130_fd_sc_hd__or2_1 _14957_ (.A(_08431_),
    .B(_08432_),
    .X(_08433_));
 sky130_vsdinv _14958_ (.A(_08433_),
    .Y(_08434_));
 sky130_fd_sc_hd__or2_1 _14959_ (.A(net286),
    .B(net318),
    .X(_08435_));
 sky130_fd_sc_hd__clkbuf_4 _14960_ (.A(net318),
    .X(_08436_));
 sky130_fd_sc_hd__nand2_1 _14961_ (.A(net286),
    .B(_08436_),
    .Y(_08437_));
 sky130_fd_sc_hd__nand2_1 _14962_ (.A(_08435_),
    .B(_08437_),
    .Y(_08438_));
 sky130_vsdinv _14963_ (.A(_08438_),
    .Y(_08439_));
 sky130_fd_sc_hd__or4_2 _14964_ (.A(_08426_),
    .B(_08430_),
    .C(_08434_),
    .D(_08439_),
    .X(_08440_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14965_ (.A(net292),
    .X(_08441_));
 sky130_fd_sc_hd__or2_1 _14966_ (.A(net186),
    .B(_08441_),
    .X(_08442_));
 sky130_fd_sc_hd__buf_1 _14967_ (.A(net186),
    .X(_08443_));
 sky130_fd_sc_hd__nand2_1 _14968_ (.A(_08443_),
    .B(_08441_),
    .Y(_08444_));
 sky130_fd_sc_hd__and2_1 _14969_ (.A(_08442_),
    .B(_08444_),
    .X(_08445_));
 sky130_fd_sc_hd__nor2_1 _14970_ (.A(net273),
    .B(net305),
    .Y(_08446_));
 sky130_fd_sc_hd__nand2_1 _14971_ (.A(net273),
    .B(net305),
    .Y(_08447_));
 sky130_fd_sc_hd__and2b_1 _14972_ (.A_N(_08446_),
    .B(_08447_),
    .X(_08448_));
 sky130_fd_sc_hd__clkbuf_2 _14973_ (.A(net294),
    .X(_08449_));
 sky130_fd_sc_hd__or2_1 _14974_ (.A(net188),
    .B(_08449_),
    .X(_08450_));
 sky130_vsdinv _14975_ (.A(_08450_),
    .Y(_08451_));
 sky130_fd_sc_hd__and2_1 _14976_ (.A(net188),
    .B(_08449_),
    .X(_08452_));
 sky130_fd_sc_hd__nor2_1 _14977_ (.A(_08451_),
    .B(_08452_),
    .Y(_08453_));
 sky130_fd_sc_hd__or2_1 _14978_ (.A(net183),
    .B(net289),
    .X(_08454_));
 sky130_fd_sc_hd__clkbuf_2 _14979_ (.A(net183),
    .X(_08455_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14980_ (.A(net289),
    .X(_08456_));
 sky130_fd_sc_hd__nand2_1 _14981_ (.A(_08455_),
    .B(_08456_),
    .Y(_08457_));
 sky130_fd_sc_hd__and2_1 _14982_ (.A(_08454_),
    .B(_08457_),
    .X(_08458_));
 sky130_fd_sc_hd__or4_1 _14983_ (.A(_08445_),
    .B(_08448_),
    .C(_08453_),
    .D(_08458_),
    .X(_08459_));
 sky130_fd_sc_hd__clkbuf_2 _14984_ (.A(net296),
    .X(_08460_));
 sky130_fd_sc_hd__clkbuf_4 _14985_ (.A(_08460_),
    .X(_08461_));
 sky130_fd_sc_hd__nor2_1 _14986_ (.A(net190),
    .B(_08461_),
    .Y(_08462_));
 sky130_fd_sc_hd__and2_1 _14987_ (.A(net190),
    .B(net296),
    .X(_08463_));
 sky130_fd_sc_hd__nor2_1 _14988_ (.A(_08462_),
    .B(_08463_),
    .Y(_08464_));
 sky130_fd_sc_hd__or2_2 _14989_ (.A(net278),
    .B(net172),
    .X(_08465_));
 sky130_fd_sc_hd__nand2_1 _14990_ (.A(_08193_),
    .B(net172),
    .Y(_08466_));
 sky130_fd_sc_hd__and2_1 _14991_ (.A(_08465_),
    .B(_08466_),
    .X(_08467_));
 sky130_vsdinv _14992_ (.A(net267),
    .Y(_08468_));
 sky130_fd_sc_hd__clkbuf_2 _14993_ (.A(net161),
    .X(_08469_));
 sky130_fd_sc_hd__inv_2 _14994_ (.A(_08469_),
    .Y(_08470_));
 sky130_fd_sc_hd__nor2_1 _14995_ (.A(_08468_),
    .B(_08470_),
    .Y(_08471_));
 sky130_fd_sc_hd__buf_2 _14996_ (.A(_08469_),
    .X(_08472_));
 sky130_fd_sc_hd__nor2_1 _14997_ (.A(_08325_),
    .B(_08472_),
    .Y(_08473_));
 sky130_fd_sc_hd__nor2_1 _14998_ (.A(_08471_),
    .B(_08473_),
    .Y(_00000_));
 sky130_fd_sc_hd__or2_1 _14999_ (.A(net187),
    .B(net293),
    .X(_08474_));
 sky130_fd_sc_hd__clkbuf_2 _15000_ (.A(net293),
    .X(_08475_));
 sky130_fd_sc_hd__nand2_1 _15001_ (.A(net187),
    .B(_08475_),
    .Y(_08476_));
 sky130_fd_sc_hd__and2_1 _15002_ (.A(_08474_),
    .B(_08476_),
    .X(_08477_));
 sky130_fd_sc_hd__nor2_1 _15003_ (.A(net287),
    .B(net319),
    .Y(_08478_));
 sky130_fd_sc_hd__clkbuf_4 _15004_ (.A(net319),
    .X(_08479_));
 sky130_fd_sc_hd__nand2_1 _15005_ (.A(net287),
    .B(_08479_),
    .Y(_08480_));
 sky130_fd_sc_hd__and2b_2 _15006_ (.A_N(_08478_),
    .B(_08480_),
    .X(_08481_));
 sky130_fd_sc_hd__clkbuf_2 _15007_ (.A(net297),
    .X(_08482_));
 sky130_fd_sc_hd__and2_1 _15008_ (.A(_08482_),
    .B(net329),
    .X(_08483_));
 sky130_fd_sc_hd__clkbuf_4 _15009_ (.A(net329),
    .X(_08484_));
 sky130_fd_sc_hd__nor2_1 _15010_ (.A(_08482_),
    .B(_08484_),
    .Y(_08485_));
 sky130_fd_sc_hd__nor2_1 _15011_ (.A(_08483_),
    .B(_08485_),
    .Y(_08486_));
 sky130_fd_sc_hd__clkbuf_4 _15012_ (.A(net322),
    .X(_08487_));
 sky130_fd_sc_hd__nand2_1 _15013_ (.A(net290),
    .B(_08487_),
    .Y(_08488_));
 sky130_fd_sc_hd__or2_1 _15014_ (.A(net290),
    .B(net322),
    .X(_08489_));
 sky130_fd_sc_hd__and2_1 _15015_ (.A(_08488_),
    .B(_08489_),
    .X(_08490_));
 sky130_fd_sc_hd__or4_1 _15016_ (.A(_08477_),
    .B(_08481_),
    .C(_08486_),
    .D(_08490_),
    .X(_08491_));
 sky130_fd_sc_hd__or4_1 _15017_ (.A(_08464_),
    .B(_08467_),
    .C(_00000_),
    .D(_08491_),
    .X(_08492_));
 sky130_fd_sc_hd__or4_1 _15018_ (.A(_08422_),
    .B(_08440_),
    .C(_08459_),
    .D(_08492_),
    .X(_08493_));
 sky130_fd_sc_hd__nor2_1 _15019_ (.A(_08406_),
    .B(_08493_),
    .Y(_00032_));
 sky130_fd_sc_hd__nor2_2 _15020_ (.A(_08183_),
    .B(_08158_),
    .Y(_08494_));
 sky130_fd_sc_hd__nand2_1 _15021_ (.A(_08311_),
    .B(alu_wait),
    .Y(_08495_));
 sky130_fd_sc_hd__clkbuf_2 _15022_ (.A(is_lui_auipc_jal),
    .X(_08496_));
 sky130_fd_sc_hd__or3_1 _15023_ (.A(_08496_),
    .B(is_slli_srli_srai),
    .C(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .X(_08497_));
 sky130_fd_sc_hd__or2b_1 _15024_ (.A(net369),
    .B_N(_08286_),
    .X(_08498_));
 sky130_fd_sc_hd__o2bb2a_1 _15025_ (.A1_N(_08180_),
    .A2_N(_08497_),
    .B1(_08498_),
    .B2(is_sb_sh_sw),
    .X(_08499_));
 sky130_fd_sc_hd__nand2_1 _15026_ (.A(_08495_),
    .B(_08499_),
    .Y(_08500_));
 sky130_fd_sc_hd__a32o_1 _15027_ (.A1(_08494_),
    .A2(_08204_),
    .A3(_08315_),
    .B1(_08500_),
    .B2(_08206_),
    .X(_00044_));
 sky130_fd_sc_hd__or3_1 _15028_ (.A(instr_slt),
    .B(instr_slti),
    .C(instr_blt),
    .X(_08501_));
 sky130_fd_sc_hd__clkbuf_1 _15029_ (.A(_08501_),
    .X(_00038_));
 sky130_fd_sc_hd__or3_1 _15030_ (.A(instr_sltu),
    .B(instr_sltiu),
    .C(instr_bltu),
    .X(_08502_));
 sky130_fd_sc_hd__clkbuf_1 _15031_ (.A(_08502_),
    .X(_00039_));
 sky130_fd_sc_hd__clkbuf_2 _15032_ (.A(_08324_),
    .X(_08503_));
 sky130_fd_sc_hd__o21a_1 _15033_ (.A1(instr_lh),
    .A2(instr_lhu),
    .B1(_08174_),
    .X(_08504_));
 sky130_fd_sc_hd__a221o_1 _15034_ (.A1(instr_sh),
    .A2(_08164_),
    .B1(_08173_),
    .B2(_08503_),
    .C1(_08504_),
    .X(_00049_));
 sky130_fd_sc_hd__clkbuf_4 _15035_ (.A(_08328_),
    .X(_08505_));
 sky130_fd_sc_hd__clkbuf_2 _15036_ (.A(_08505_),
    .X(_08506_));
 sky130_fd_sc_hd__and3_1 _15037_ (.A(_08163_),
    .B(_08506_),
    .C(_08154_),
    .X(_08507_));
 sky130_fd_sc_hd__buf_1 _15038_ (.A(_08507_),
    .X(net193));
 sky130_fd_sc_hd__buf_2 _15039_ (.A(\mem_wordsize[1] ),
    .X(_08508_));
 sky130_fd_sc_hd__clkbuf_2 _15040_ (.A(_08508_),
    .X(_08509_));
 sky130_fd_sc_hd__clkbuf_2 _15041_ (.A(_08509_),
    .X(_08510_));
 sky130_fd_sc_hd__buf_2 _15042_ (.A(_08510_),
    .X(_08511_));
 sky130_fd_sc_hd__o21a_1 _15043_ (.A1(instr_lb),
    .A2(instr_lbu),
    .B1(_08174_),
    .X(_08512_));
 sky130_fd_sc_hd__a221o_1 _15044_ (.A1(instr_sb),
    .A2(_08164_),
    .B1(_08173_),
    .B2(_08511_),
    .C1(_08512_),
    .X(_00048_));
 sky130_vsdinv _15045_ (.A(\cpu_state[2] ),
    .Y(_08513_));
 sky130_fd_sc_hd__or2_1 _15046_ (.A(_08513_),
    .B(_08224_),
    .X(_08514_));
 sky130_fd_sc_hd__nor2_1 _15047_ (.A(_08497_),
    .B(_08514_),
    .Y(_08515_));
 sky130_fd_sc_hd__and2_1 _15048_ (.A(_08282_),
    .B(_08320_),
    .X(_08516_));
 sky130_fd_sc_hd__o211a_1 _15049_ (.A1(_08515_),
    .A2(_08516_),
    .B1(_08206_),
    .C1(_08226_),
    .X(_00043_));
 sky130_fd_sc_hd__buf_2 _15050_ (.A(_08287_),
    .X(_08517_));
 sky130_fd_sc_hd__clkbuf_2 _15051_ (.A(_08517_),
    .X(_08518_));
 sky130_fd_sc_hd__buf_2 _15052_ (.A(is_sb_sh_sw),
    .X(_08519_));
 sky130_fd_sc_hd__a32o_1 _15053_ (.A1(_08518_),
    .A2(_08519_),
    .A3(_08206_),
    .B1(_08229_),
    .B2(\cpu_state[5] ),
    .X(_00045_));
 sky130_fd_sc_hd__clkbuf_4 _15054_ (.A(_08183_),
    .X(_08520_));
 sky130_fd_sc_hd__buf_2 _15055_ (.A(_08520_),
    .X(_08521_));
 sky130_fd_sc_hd__clkbuf_2 _15056_ (.A(mem_do_rinst),
    .X(_08522_));
 sky130_fd_sc_hd__or2_1 _15057_ (.A(_08522_),
    .B(_08153_),
    .X(_08523_));
 sky130_fd_sc_hd__o21ai_2 _15058_ (.A1(_08151_),
    .A2(_08523_),
    .B1(_08154_),
    .Y(_08524_));
 sky130_fd_sc_hd__buf_2 _15059_ (.A(_08524_),
    .X(_08525_));
 sky130_fd_sc_hd__nor2_1 _15060_ (.A(_08521_),
    .B(_08525_),
    .Y(net160));
 sky130_fd_sc_hd__buf_2 _15061_ (.A(_08290_),
    .X(_08526_));
 sky130_fd_sc_hd__clkbuf_4 _15062_ (.A(_08526_),
    .X(_08527_));
 sky130_fd_sc_hd__mux2_1 _15063_ (.A0(instr_bge),
    .A1(is_slti_blt_slt),
    .S(alu_lts),
    .X(_08528_));
 sky130_vsdinv _15064_ (.A(alu_eq),
    .Y(_08529_));
 sky130_fd_sc_hd__and2b_1 _15065_ (.A_N(alu_ltu),
    .B(instr_bgeu),
    .X(_08530_));
 sky130_fd_sc_hd__a221o_1 _15066_ (.A1(instr_bne),
    .A2(_08529_),
    .B1(is_sltiu_bltu_sltu),
    .B2(alu_ltu),
    .C1(_08530_),
    .X(_08531_));
 sky130_fd_sc_hd__or4_1 _15067_ (.A(instr_bgeu),
    .B(instr_bge),
    .C(_08529_),
    .D(is_sltiu_bltu_sltu),
    .X(_08532_));
 sky130_fd_sc_hd__or3_1 _15068_ (.A(instr_bne),
    .B(is_slti_blt_slt),
    .C(_08532_),
    .X(_08533_));
 sky130_fd_sc_hd__or3b_4 _15069_ (.A(_08528_),
    .B(_08531_),
    .C_N(_08533_),
    .X(_08534_));
 sky130_fd_sc_hd__nand3_1 _15070_ (.A(_08522_),
    .B(_08328_),
    .C(_08157_),
    .Y(_08535_));
 sky130_fd_sc_hd__clkbuf_4 _15071_ (.A(_08535_),
    .X(_08536_));
 sky130_fd_sc_hd__a31o_1 _15072_ (.A1(_08527_),
    .A2(_08315_),
    .A3(_08534_),
    .B1(_08536_),
    .X(_08537_));
 sky130_fd_sc_hd__nand2_1 _15073_ (.A(_08292_),
    .B(_08537_),
    .Y(_00035_));
 sky130_fd_sc_hd__or2_2 _15074_ (.A(\cpu_state[2] ),
    .B(_08286_),
    .X(_08538_));
 sky130_fd_sc_hd__or2_1 _15075_ (.A(\cpu_state[4] ),
    .B(_08538_),
    .X(_08539_));
 sky130_fd_sc_hd__or2_1 _15076_ (.A(\cpu_state[6] ),
    .B(_08539_),
    .X(_08540_));
 sky130_fd_sc_hd__clkbuf_2 _15077_ (.A(_08540_),
    .X(_08541_));
 sky130_fd_sc_hd__clkbuf_2 _15078_ (.A(_08541_),
    .X(_08542_));
 sky130_fd_sc_hd__mux2_2 _15079_ (.A0(\decoded_rs1[4] ),
    .A1(\decoded_imm_uj[4] ),
    .S(_08285_),
    .X(_08543_));
 sky130_fd_sc_hd__buf_2 _15080_ (.A(_08543_),
    .X(_08544_));
 sky130_fd_sc_hd__clkbuf_4 _15081_ (.A(_08544_),
    .X(_08545_));
 sky130_fd_sc_hd__buf_2 _15082_ (.A(\decoded_imm_uj[1] ),
    .X(_08546_));
 sky130_vsdinv _15083_ (.A(_08546_),
    .Y(_08547_));
 sky130_fd_sc_hd__nand2_1 _15084_ (.A(_08284_),
    .B(_08547_),
    .Y(_08548_));
 sky130_fd_sc_hd__o21a_2 _15085_ (.A1(_08284_),
    .A2(\decoded_rs1[1] ),
    .B1(_08548_),
    .X(_08549_));
 sky130_fd_sc_hd__clkbuf_4 _15086_ (.A(_08549_),
    .X(_08550_));
 sky130_fd_sc_hd__clkbuf_2 _15087_ (.A(_08550_),
    .X(_08551_));
 sky130_fd_sc_hd__buf_2 _15088_ (.A(_08551_),
    .X(_08552_));
 sky130_fd_sc_hd__buf_2 _15089_ (.A(_08552_),
    .X(_08553_));
 sky130_fd_sc_hd__clkbuf_4 _15090_ (.A(\decoded_imm_uj[11] ),
    .X(_08554_));
 sky130_fd_sc_hd__or2b_1 _15091_ (.A(_08554_),
    .B_N(\cpu_state[3] ),
    .X(_08555_));
 sky130_fd_sc_hd__o21a_4 _15092_ (.A1(\cpu_state[3] ),
    .A2(\decoded_rs1[0] ),
    .B1(_08555_),
    .X(_08556_));
 sky130_fd_sc_hd__clkbuf_2 _15093_ (.A(_08556_),
    .X(_08557_));
 sky130_fd_sc_hd__clkbuf_2 _15094_ (.A(_08557_),
    .X(_08558_));
 sky130_fd_sc_hd__buf_4 _15095_ (.A(_08558_),
    .X(_08559_));
 sky130_fd_sc_hd__buf_2 _15096_ (.A(_08559_),
    .X(_08560_));
 sky130_fd_sc_hd__clkbuf_4 _15097_ (.A(_08560_),
    .X(_08561_));
 sky130_fd_sc_hd__mux2_1 _15098_ (.A0(\cpuregs[18][0] ),
    .A1(\cpuregs[19][0] ),
    .S(_08561_),
    .X(_08562_));
 sky130_fd_sc_hd__o21ai_1 _15099_ (.A1(_08286_),
    .A2(\decoded_rs1[0] ),
    .B1(_08555_),
    .Y(_08563_));
 sky130_fd_sc_hd__clkbuf_2 _15100_ (.A(_08563_),
    .X(_08564_));
 sky130_fd_sc_hd__buf_2 _15101_ (.A(_08564_),
    .X(_08565_));
 sky130_fd_sc_hd__o21ai_2 _15102_ (.A1(_08284_),
    .A2(\decoded_rs1[1] ),
    .B1(_08548_),
    .Y(_08566_));
 sky130_fd_sc_hd__clkbuf_2 _15103_ (.A(_08566_),
    .X(_08567_));
 sky130_fd_sc_hd__clkbuf_4 _15104_ (.A(_08567_),
    .X(_08568_));
 sky130_fd_sc_hd__clkbuf_4 _15105_ (.A(_08568_),
    .X(_08569_));
 sky130_fd_sc_hd__clkbuf_2 _15106_ (.A(_08569_),
    .X(_08570_));
 sky130_fd_sc_hd__buf_2 _15107_ (.A(_08557_),
    .X(_08571_));
 sky130_fd_sc_hd__buf_2 _15108_ (.A(_08571_),
    .X(_08572_));
 sky130_fd_sc_hd__clkbuf_4 _15109_ (.A(_08572_),
    .X(_08573_));
 sky130_fd_sc_hd__buf_2 _15110_ (.A(_08573_),
    .X(_08574_));
 sky130_fd_sc_hd__or2_1 _15111_ (.A(\cpuregs[16][0] ),
    .B(_08574_),
    .X(_08575_));
 sky130_fd_sc_hd__o211a_1 _15112_ (.A1(\cpuregs[17][0] ),
    .A2(_08565_),
    .B1(_08570_),
    .C1(_08575_),
    .X(_08576_));
 sky130_fd_sc_hd__a21oi_1 _15113_ (.A1(_08553_),
    .A2(_08562_),
    .B1(_08576_),
    .Y(_08577_));
 sky130_fd_sc_hd__or2b_1 _15114_ (.A(\decoded_imm_uj[2] ),
    .B_N(_08284_),
    .X(_08578_));
 sky130_fd_sc_hd__o21ai_4 _15115_ (.A1(_08285_),
    .A2(\decoded_rs1[2] ),
    .B1(_08578_),
    .Y(_08579_));
 sky130_fd_sc_hd__clkbuf_2 _15116_ (.A(_08579_),
    .X(_08580_));
 sky130_fd_sc_hd__clkbuf_4 _15117_ (.A(_08580_),
    .X(_08581_));
 sky130_fd_sc_hd__clkbuf_4 _15118_ (.A(_08571_),
    .X(_08582_));
 sky130_fd_sc_hd__mux2_1 _15119_ (.A0(\cpuregs[10][0] ),
    .A1(\cpuregs[11][0] ),
    .S(_08582_),
    .X(_08583_));
 sky130_fd_sc_hd__mux2_1 _15120_ (.A0(\cpuregs[8][0] ),
    .A1(\cpuregs[9][0] ),
    .S(_08582_),
    .X(_08584_));
 sky130_fd_sc_hd__buf_2 _15121_ (.A(_08566_),
    .X(_08585_));
 sky130_fd_sc_hd__buf_4 _15122_ (.A(_08585_),
    .X(_08586_));
 sky130_fd_sc_hd__mux2_1 _15123_ (.A0(_08583_),
    .A1(_08584_),
    .S(_08586_),
    .X(_08587_));
 sky130_fd_sc_hd__buf_1 _15124_ (.A(_08549_),
    .X(_08588_));
 sky130_fd_sc_hd__buf_2 _15125_ (.A(_08588_),
    .X(_08589_));
 sky130_fd_sc_hd__buf_2 _15126_ (.A(_08558_),
    .X(_08590_));
 sky130_fd_sc_hd__mux2_1 _15127_ (.A0(\cpuregs[12][0] ),
    .A1(\cpuregs[13][0] ),
    .S(_08590_),
    .X(_08591_));
 sky130_fd_sc_hd__clkbuf_2 _15128_ (.A(_08566_),
    .X(_08592_));
 sky130_fd_sc_hd__clkbuf_4 _15129_ (.A(_08592_),
    .X(_08593_));
 sky130_fd_sc_hd__clkbuf_2 _15130_ (.A(_08556_),
    .X(_08594_));
 sky130_fd_sc_hd__buf_4 _15131_ (.A(_08594_),
    .X(_08595_));
 sky130_fd_sc_hd__mux2_1 _15132_ (.A0(\cpuregs[14][0] ),
    .A1(\cpuregs[15][0] ),
    .S(_08595_),
    .X(_08596_));
 sky130_fd_sc_hd__or2_1 _15133_ (.A(_08593_),
    .B(_08596_),
    .X(_08597_));
 sky130_fd_sc_hd__o21a_2 _15134_ (.A1(_08285_),
    .A2(\decoded_rs1[2] ),
    .B1(_08578_),
    .X(_08598_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15135_ (.A(_08598_),
    .X(_08599_));
 sky130_fd_sc_hd__clkbuf_4 _15136_ (.A(_08599_),
    .X(_08600_));
 sky130_fd_sc_hd__o211a_1 _15137_ (.A1(_08589_),
    .A2(_08591_),
    .B1(_08597_),
    .C1(_08600_),
    .X(_08601_));
 sky130_fd_sc_hd__or2b_1 _15138_ (.A(\decoded_imm_uj[3] ),
    .B_N(_08284_),
    .X(_08602_));
 sky130_fd_sc_hd__o21ai_2 _15139_ (.A1(_08285_),
    .A2(\decoded_rs1[3] ),
    .B1(_08602_),
    .Y(_08603_));
 sky130_fd_sc_hd__buf_2 _15140_ (.A(_08603_),
    .X(_08604_));
 sky130_fd_sc_hd__buf_2 _15141_ (.A(_08604_),
    .X(_08605_));
 sky130_fd_sc_hd__a211o_1 _15142_ (.A1(_08581_),
    .A2(_08587_),
    .B1(_08601_),
    .C1(_08605_),
    .X(_08606_));
 sky130_fd_sc_hd__buf_2 _15143_ (.A(_08579_),
    .X(_08607_));
 sky130_fd_sc_hd__clkbuf_4 _15144_ (.A(_08607_),
    .X(_08608_));
 sky130_fd_sc_hd__clkbuf_2 _15145_ (.A(_08556_),
    .X(_08609_));
 sky130_fd_sc_hd__clkbuf_4 _15146_ (.A(_08609_),
    .X(_08610_));
 sky130_fd_sc_hd__mux2_1 _15147_ (.A0(\cpuregs[2][0] ),
    .A1(\cpuregs[3][0] ),
    .S(_08610_),
    .X(_08611_));
 sky130_fd_sc_hd__mux2_1 _15148_ (.A0(\cpuregs[0][0] ),
    .A1(\cpuregs[1][0] ),
    .S(_08610_),
    .X(_08612_));
 sky130_fd_sc_hd__clkbuf_4 _15149_ (.A(_08567_),
    .X(_08613_));
 sky130_fd_sc_hd__mux2_1 _15150_ (.A0(_08611_),
    .A1(_08612_),
    .S(_08613_),
    .X(_08614_));
 sky130_fd_sc_hd__o21a_1 _15151_ (.A1(_08285_),
    .A2(\decoded_rs1[3] ),
    .B1(_08602_),
    .X(_08615_));
 sky130_fd_sc_hd__buf_2 _15152_ (.A(_08615_),
    .X(_08616_));
 sky130_fd_sc_hd__buf_2 _15153_ (.A(_08616_),
    .X(_08617_));
 sky130_fd_sc_hd__buf_4 _15154_ (.A(_08558_),
    .X(_08618_));
 sky130_fd_sc_hd__mux2_1 _15155_ (.A0(\cpuregs[4][0] ),
    .A1(\cpuregs[5][0] ),
    .S(_08618_),
    .X(_08619_));
 sky130_fd_sc_hd__buf_2 _15156_ (.A(_08599_),
    .X(_08620_));
 sky130_fd_sc_hd__clkbuf_4 _15157_ (.A(_08594_),
    .X(_08621_));
 sky130_fd_sc_hd__mux2_1 _15158_ (.A0(\cpuregs[6][0] ),
    .A1(\cpuregs[7][0] ),
    .S(_08621_),
    .X(_08622_));
 sky130_fd_sc_hd__or2_1 _15159_ (.A(_08568_),
    .B(_08622_),
    .X(_08623_));
 sky130_fd_sc_hd__o211a_1 _15160_ (.A1(_08589_),
    .A2(_08619_),
    .B1(_08620_),
    .C1(_08623_),
    .X(_08624_));
 sky130_fd_sc_hd__a211o_1 _15161_ (.A1(_08608_),
    .A2(_08614_),
    .B1(_08617_),
    .C1(_08624_),
    .X(_08625_));
 sky130_fd_sc_hd__buf_2 _15162_ (.A(_08543_),
    .X(_08626_));
 sky130_fd_sc_hd__clkbuf_4 _15163_ (.A(_08626_),
    .X(_08627_));
 sky130_fd_sc_hd__a21oi_2 _15164_ (.A1(_08606_),
    .A2(_08625_),
    .B1(_08627_),
    .Y(_08628_));
 sky130_fd_sc_hd__buf_2 _15165_ (.A(_08560_),
    .X(_08629_));
 sky130_fd_sc_hd__clkbuf_2 _15166_ (.A(_08549_),
    .X(_08630_));
 sky130_fd_sc_hd__or4_1 _15167_ (.A(_08630_),
    .B(_08598_),
    .C(_08615_),
    .D(_08543_),
    .X(_08631_));
 sky130_fd_sc_hd__nor2_1 _15168_ (.A(_08629_),
    .B(_08631_),
    .Y(_08632_));
 sky130_fd_sc_hd__clkbuf_2 _15169_ (.A(_08632_),
    .X(_08633_));
 sky130_fd_sc_hd__clkbuf_4 _15170_ (.A(_08633_),
    .X(_08634_));
 sky130_fd_sc_hd__a211o_4 _15171_ (.A1(_08545_),
    .A2(_08577_),
    .B1(_08628_),
    .C1(_08634_),
    .X(_08635_));
 sky130_fd_sc_hd__o21ba_1 _15172_ (.A1(instr_getq),
    .A2(instr_setq),
    .B1_N(_08635_),
    .X(_08636_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15173_ (.A(instr_maskirq),
    .X(_08637_));
 sky130_fd_sc_hd__clkbuf_2 _15174_ (.A(_08637_),
    .X(_08638_));
 sky130_fd_sc_hd__clkbuf_2 _15175_ (.A(_08638_),
    .X(_08639_));
 sky130_fd_sc_hd__clkbuf_2 _15176_ (.A(instr_timer),
    .X(_08640_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15177_ (.A(_08640_),
    .X(_08641_));
 sky130_fd_sc_hd__clkbuf_2 _15178_ (.A(_08641_),
    .X(_08642_));
 sky130_fd_sc_hd__clkbuf_2 _15179_ (.A(_08642_),
    .X(_08643_));
 sky130_fd_sc_hd__nor3b_1 _15180_ (.A(_08640_),
    .B(instr_maskirq),
    .C_N(_08221_),
    .Y(_08644_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15181_ (.A(_08644_),
    .X(_08645_));
 sky130_fd_sc_hd__clkbuf_2 _15182_ (.A(_08645_),
    .X(_08646_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15183_ (.A(_08646_),
    .X(_08647_));
 sky130_fd_sc_hd__a221o_1 _15184_ (.A1(\irq_mask[0] ),
    .A2(_08639_),
    .B1(\timer[0] ),
    .B2(_08643_),
    .C1(_08647_),
    .X(_08648_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15185_ (.A(_08222_),
    .X(_08649_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15186_ (.A(_08649_),
    .X(_08650_));
 sky130_fd_sc_hd__clkbuf_2 _15187_ (.A(instr_rdcycleh),
    .X(_08651_));
 sky130_fd_sc_hd__clkbuf_2 _15188_ (.A(_08651_),
    .X(_08652_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15189_ (.A(net373),
    .X(_08653_));
 sky130_fd_sc_hd__buf_2 _15190_ (.A(_08653_),
    .X(_08654_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15191_ (.A(\count_cycle[0] ),
    .X(_08655_));
 sky130_fd_sc_hd__clkbuf_2 _15192_ (.A(instr_rdinstr),
    .X(_08656_));
 sky130_fd_sc_hd__clkbuf_2 _15193_ (.A(instr_rdinstrh),
    .X(_08657_));
 sky130_fd_sc_hd__clkbuf_2 _15194_ (.A(_08657_),
    .X(_08658_));
 sky130_fd_sc_hd__a22o_1 _15195_ (.A1(\count_instr[0] ),
    .A2(_08656_),
    .B1(_08658_),
    .B2(\count_instr[32] ),
    .X(_08659_));
 sky130_fd_sc_hd__a221o_1 _15196_ (.A1(_08652_),
    .A2(\count_cycle[32] ),
    .B1(_08654_),
    .B2(_08655_),
    .C1(_08659_),
    .X(_08660_));
 sky130_fd_sc_hd__or2_1 _15197_ (.A(_08650_),
    .B(_08660_),
    .X(_08661_));
 sky130_fd_sc_hd__o211a_1 _15198_ (.A1(_08636_),
    .A2(_08648_),
    .B1(_08661_),
    .C1(_08181_),
    .X(_08662_));
 sky130_fd_sc_hd__nor2_1 _15199_ (.A(\cpu_state[6] ),
    .B(_08539_),
    .Y(_08663_));
 sky130_fd_sc_hd__clkbuf_2 _15200_ (.A(_08663_),
    .X(_08664_));
 sky130_fd_sc_hd__clkbuf_2 _15201_ (.A(_08664_),
    .X(_08665_));
 sky130_fd_sc_hd__clkbuf_2 _15202_ (.A(_08665_),
    .X(_08666_));
 sky130_fd_sc_hd__clkbuf_2 _15203_ (.A(\reg_next_pc[0] ),
    .X(_08667_));
 sky130_fd_sc_hd__clkbuf_2 _15204_ (.A(\decoded_imm[0] ),
    .X(_08668_));
 sky130_fd_sc_hd__o21ai_1 _15205_ (.A1(_08667_),
    .A2(_08668_),
    .B1(_08312_),
    .Y(_08669_));
 sky130_fd_sc_hd__a21oi_1 _15206_ (.A1(_08667_),
    .A2(_08668_),
    .B1(_08669_),
    .Y(_08670_));
 sky130_fd_sc_hd__clkbuf_2 _15207_ (.A(_08152_),
    .X(_08671_));
 sky130_vsdinv _15208_ (.A(_08193_),
    .Y(_08672_));
 sky130_fd_sc_hd__nor2_2 _15209_ (.A(\mem_wordsize[2] ),
    .B(\mem_wordsize[1] ),
    .Y(_08673_));
 sky130_fd_sc_hd__nor2_1 _15210_ (.A(_08672_),
    .B(_08673_),
    .Y(_08674_));
 sky130_fd_sc_hd__o21a_1 _15211_ (.A1(\mem_wordsize[2] ),
    .A2(_08468_),
    .B1(_08674_),
    .X(_08675_));
 sky130_fd_sc_hd__nand2_1 _15212_ (.A(\mem_wordsize[2] ),
    .B(_08193_),
    .Y(_08676_));
 sky130_fd_sc_hd__nand2b_4 _15213_ (.A_N(\mem_wordsize[2] ),
    .B(_08508_),
    .Y(_08677_));
 sky130_fd_sc_hd__a22o_1 _15214_ (.A1(_08468_),
    .A2(_08672_),
    .B1(_08676_),
    .B2(_08677_),
    .X(_08678_));
 sky130_fd_sc_hd__buf_2 _15215_ (.A(_08193_),
    .X(_08679_));
 sky130_fd_sc_hd__o211a_1 _15216_ (.A1(_08679_),
    .A2(net63),
    .B1(_08508_),
    .C1(_08191_),
    .X(_08680_));
 sky130_fd_sc_hd__o21a_1 _15217_ (.A1(_08672_),
    .A2(net49),
    .B1(_08680_),
    .X(_08681_));
 sky130_fd_sc_hd__a221o_1 _15218_ (.A1(net40),
    .A2(_08675_),
    .B1(_08678_),
    .B2(net33),
    .C1(_08681_),
    .X(_08682_));
 sky130_fd_sc_hd__clkbuf_2 _15219_ (.A(\genblk1.pcpi_mul.shift_out ),
    .X(_08683_));
 sky130_fd_sc_hd__mux2_2 _15220_ (.A0(\genblk1.pcpi_mul.rd[0] ),
    .A1(\genblk1.pcpi_mul.rd[32] ),
    .S(_08683_),
    .X(_08684_));
 sky130_fd_sc_hd__clkbuf_2 _15221_ (.A(_08286_),
    .X(_08685_));
 sky130_fd_sc_hd__a22o_1 _15222_ (.A1(_08671_),
    .A2(_08682_),
    .B1(_08684_),
    .B2(_08685_),
    .X(_08686_));
 sky130_fd_sc_hd__or3_1 _15223_ (.A(_08666_),
    .B(_08670_),
    .C(_08686_),
    .X(_08687_));
 sky130_fd_sc_hd__o22a_1 _15224_ (.A1(\irq_pending[0] ),
    .A2(_08542_),
    .B1(_08662_),
    .B2(_08687_),
    .X(_14572_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15225_ (.A(_08221_),
    .X(_08688_));
 sky130_fd_sc_hd__clkbuf_2 _15226_ (.A(_08688_),
    .X(_08689_));
 sky130_fd_sc_hd__clkbuf_2 _15227_ (.A(_08689_),
    .X(_08690_));
 sky130_fd_sc_hd__clkbuf_4 _15228_ (.A(_08543_),
    .X(_08691_));
 sky130_fd_sc_hd__buf_2 _15229_ (.A(_08691_),
    .X(_08692_));
 sky130_fd_sc_hd__buf_2 _15230_ (.A(_08552_),
    .X(_08693_));
 sky130_fd_sc_hd__clkbuf_2 _15231_ (.A(_08556_),
    .X(_08694_));
 sky130_fd_sc_hd__buf_2 _15232_ (.A(_08694_),
    .X(_08695_));
 sky130_fd_sc_hd__clkbuf_4 _15233_ (.A(_08695_),
    .X(_08696_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15234_ (.A(_08696_),
    .X(_08697_));
 sky130_fd_sc_hd__buf_2 _15235_ (.A(_08697_),
    .X(_08698_));
 sky130_fd_sc_hd__mux2_1 _15236_ (.A0(\cpuregs[18][1] ),
    .A1(\cpuregs[19][1] ),
    .S(_08698_),
    .X(_08699_));
 sky130_fd_sc_hd__clkbuf_2 _15237_ (.A(_08564_),
    .X(_08700_));
 sky130_fd_sc_hd__clkbuf_2 _15238_ (.A(_08569_),
    .X(_08701_));
 sky130_fd_sc_hd__buf_2 _15239_ (.A(_08701_),
    .X(_08702_));
 sky130_fd_sc_hd__or2_1 _15240_ (.A(\cpuregs[16][1] ),
    .B(_08698_),
    .X(_08703_));
 sky130_fd_sc_hd__o211a_1 _15241_ (.A1(\cpuregs[17][1] ),
    .A2(_08700_),
    .B1(_08702_),
    .C1(_08703_),
    .X(_08704_));
 sky130_fd_sc_hd__a21oi_1 _15242_ (.A1(_08693_),
    .A2(_08699_),
    .B1(_08704_),
    .Y(_08705_));
 sky130_fd_sc_hd__clkbuf_2 _15243_ (.A(_08579_),
    .X(_08706_));
 sky130_fd_sc_hd__clkbuf_4 _15244_ (.A(_08706_),
    .X(_08707_));
 sky130_fd_sc_hd__buf_2 _15245_ (.A(_08707_),
    .X(_08708_));
 sky130_fd_sc_hd__clkbuf_4 _15246_ (.A(_08571_),
    .X(_08709_));
 sky130_fd_sc_hd__buf_2 _15247_ (.A(_08709_),
    .X(_08710_));
 sky130_fd_sc_hd__mux2_1 _15248_ (.A0(\cpuregs[8][1] ),
    .A1(\cpuregs[9][1] ),
    .S(_08710_),
    .X(_08711_));
 sky130_fd_sc_hd__mux2_1 _15249_ (.A0(\cpuregs[10][1] ),
    .A1(\cpuregs[11][1] ),
    .S(_08710_),
    .X(_08712_));
 sky130_fd_sc_hd__clkbuf_2 _15250_ (.A(_08549_),
    .X(_08713_));
 sky130_fd_sc_hd__clkbuf_4 _15251_ (.A(_08713_),
    .X(_08714_));
 sky130_fd_sc_hd__mux2_1 _15252_ (.A0(_08711_),
    .A1(_08712_),
    .S(_08714_),
    .X(_08715_));
 sky130_fd_sc_hd__clkbuf_4 _15253_ (.A(_08589_),
    .X(_08716_));
 sky130_fd_sc_hd__clkbuf_4 _15254_ (.A(_08694_),
    .X(_08717_));
 sky130_fd_sc_hd__clkbuf_4 _15255_ (.A(_08717_),
    .X(_08718_));
 sky130_fd_sc_hd__clkbuf_4 _15256_ (.A(_08718_),
    .X(_08719_));
 sky130_fd_sc_hd__mux2_1 _15257_ (.A0(\cpuregs[12][1] ),
    .A1(\cpuregs[13][1] ),
    .S(_08719_),
    .X(_08720_));
 sky130_fd_sc_hd__buf_2 _15258_ (.A(_08593_),
    .X(_08721_));
 sky130_fd_sc_hd__mux2_1 _15259_ (.A0(\cpuregs[14][1] ),
    .A1(\cpuregs[15][1] ),
    .S(_08718_),
    .X(_08722_));
 sky130_fd_sc_hd__or2_1 _15260_ (.A(_08721_),
    .B(_08722_),
    .X(_08723_));
 sky130_fd_sc_hd__buf_2 _15261_ (.A(_08600_),
    .X(_08724_));
 sky130_fd_sc_hd__o211a_1 _15262_ (.A1(_08716_),
    .A2(_08720_),
    .B1(_08723_),
    .C1(_08724_),
    .X(_08725_));
 sky130_fd_sc_hd__clkbuf_4 _15263_ (.A(_08604_),
    .X(_08726_));
 sky130_fd_sc_hd__a211o_1 _15264_ (.A1(_08708_),
    .A2(_08715_),
    .B1(_08725_),
    .C1(_08726_),
    .X(_08727_));
 sky130_fd_sc_hd__mux2_1 _15265_ (.A0(\cpuregs[6][1] ),
    .A1(\cpuregs[7][1] ),
    .S(_08710_),
    .X(_08728_));
 sky130_fd_sc_hd__mux2_1 _15266_ (.A0(\cpuregs[4][1] ),
    .A1(\cpuregs[5][1] ),
    .S(_08710_),
    .X(_08729_));
 sky130_fd_sc_hd__buf_2 _15267_ (.A(_08592_),
    .X(_08730_));
 sky130_fd_sc_hd__buf_2 _15268_ (.A(_08730_),
    .X(_08731_));
 sky130_fd_sc_hd__clkbuf_4 _15269_ (.A(_08731_),
    .X(_08732_));
 sky130_fd_sc_hd__mux2_1 _15270_ (.A0(_08728_),
    .A1(_08729_),
    .S(_08732_),
    .X(_08733_));
 sky130_fd_sc_hd__mux2_1 _15271_ (.A0(\cpuregs[0][1] ),
    .A1(\cpuregs[1][1] ),
    .S(_08719_),
    .X(_08734_));
 sky130_fd_sc_hd__buf_2 _15272_ (.A(_08592_),
    .X(_08735_));
 sky130_fd_sc_hd__clkbuf_2 _15273_ (.A(_08735_),
    .X(_08736_));
 sky130_fd_sc_hd__mux2_1 _15274_ (.A0(\cpuregs[2][1] ),
    .A1(\cpuregs[3][1] ),
    .S(_08618_),
    .X(_08737_));
 sky130_fd_sc_hd__or2_1 _15275_ (.A(_08736_),
    .B(_08737_),
    .X(_08738_));
 sky130_fd_sc_hd__o211a_1 _15276_ (.A1(_08716_),
    .A2(_08734_),
    .B1(_08738_),
    .C1(_08581_),
    .X(_08739_));
 sky130_fd_sc_hd__clkbuf_4 _15277_ (.A(_08616_),
    .X(_08740_));
 sky130_fd_sc_hd__a211o_1 _15278_ (.A1(_08724_),
    .A2(_08733_),
    .B1(_08739_),
    .C1(_08740_),
    .X(_08741_));
 sky130_fd_sc_hd__a21oi_1 _15279_ (.A1(_08727_),
    .A2(_08741_),
    .B1(_08692_),
    .Y(_08742_));
 sky130_fd_sc_hd__clkbuf_4 _15280_ (.A(_08633_),
    .X(_08743_));
 sky130_fd_sc_hd__a211o_4 _15281_ (.A1(_08692_),
    .A2(_08705_),
    .B1(_08742_),
    .C1(_08743_),
    .X(_08744_));
 sky130_fd_sc_hd__nor2_1 _15282_ (.A(_08690_),
    .B(_08744_),
    .Y(_08745_));
 sky130_fd_sc_hd__a221o_1 _15283_ (.A1(_08281_),
    .A2(_08639_),
    .B1(\timer[1] ),
    .B2(_08643_),
    .C1(_08647_),
    .X(_08746_));
 sky130_fd_sc_hd__clkbuf_2 _15284_ (.A(_08653_),
    .X(_08747_));
 sky130_fd_sc_hd__clkbuf_2 _15285_ (.A(_08747_),
    .X(_08748_));
 sky130_fd_sc_hd__buf_2 _15286_ (.A(_08656_),
    .X(_08749_));
 sky130_fd_sc_hd__a22o_1 _15287_ (.A1(\count_instr[33] ),
    .A2(_08658_),
    .B1(_08652_),
    .B2(\count_cycle[33] ),
    .X(_08750_));
 sky130_fd_sc_hd__a21o_1 _15288_ (.A1(\count_instr[1] ),
    .A2(_08749_),
    .B1(_08750_),
    .X(_08751_));
 sky130_fd_sc_hd__clkbuf_2 _15289_ (.A(_08222_),
    .X(_08752_));
 sky130_fd_sc_hd__clkbuf_2 _15290_ (.A(_08752_),
    .X(_08753_));
 sky130_fd_sc_hd__a211o_1 _15291_ (.A1(\count_cycle[1] ),
    .A2(_08748_),
    .B1(_08751_),
    .C1(_08753_),
    .X(_08754_));
 sky130_fd_sc_hd__o211a_1 _15292_ (.A1(_08745_),
    .A2(_08746_),
    .B1(_08754_),
    .C1(_08181_),
    .X(_08755_));
 sky130_fd_sc_hd__clkbuf_2 _15293_ (.A(_08675_),
    .X(_08756_));
 sky130_fd_sc_hd__buf_2 _15294_ (.A(_08678_),
    .X(net194));
 sky130_fd_sc_hd__buf_2 _15295_ (.A(_08672_),
    .X(_08757_));
 sky130_fd_sc_hd__buf_2 _15296_ (.A(_08679_),
    .X(_08758_));
 sky130_fd_sc_hd__o211a_1 _15297_ (.A1(_08758_),
    .A2(net64),
    .B1(_08509_),
    .C1(_08326_),
    .X(_08759_));
 sky130_fd_sc_hd__o21a_1 _15298_ (.A1(_08757_),
    .A2(net50),
    .B1(_08759_),
    .X(_08760_));
 sky130_fd_sc_hd__a221o_1 _15299_ (.A1(net41),
    .A2(_08756_),
    .B1(net194),
    .B2(net44),
    .C1(_08760_),
    .X(_08761_));
 sky130_fd_sc_hd__clkbuf_2 _15300_ (.A(\decoded_imm[1] ),
    .X(_08762_));
 sky130_fd_sc_hd__nand2_1 _15301_ (.A(_08184_),
    .B(_08762_),
    .Y(_08763_));
 sky130_fd_sc_hd__or2_1 _15302_ (.A(\reg_pc[1] ),
    .B(_08762_),
    .X(_08764_));
 sky130_fd_sc_hd__and4_1 _15303_ (.A(_08667_),
    .B(\decoded_imm[0] ),
    .C(_08763_),
    .D(_08764_),
    .X(_08765_));
 sky130_vsdinv _15304_ (.A(_08765_),
    .Y(_08766_));
 sky130_fd_sc_hd__a22o_1 _15305_ (.A1(_08667_),
    .A2(\decoded_imm[0] ),
    .B1(_08763_),
    .B2(_08764_),
    .X(_08767_));
 sky130_fd_sc_hd__buf_2 _15306_ (.A(\genblk1.pcpi_mul.shift_out ),
    .X(_08768_));
 sky130_fd_sc_hd__buf_2 _15307_ (.A(_08768_),
    .X(_08769_));
 sky130_fd_sc_hd__mux2_2 _15308_ (.A0(\genblk1.pcpi_mul.rd[1] ),
    .A1(\genblk1.pcpi_mul.rd[33] ),
    .S(_08769_),
    .X(_08770_));
 sky130_fd_sc_hd__buf_2 _15309_ (.A(_08287_),
    .X(_08771_));
 sky130_fd_sc_hd__a32o_1 _15310_ (.A1(_08312_),
    .A2(_08766_),
    .A3(_08767_),
    .B1(_08770_),
    .B2(_08771_),
    .X(_08772_));
 sky130_fd_sc_hd__clkbuf_2 _15311_ (.A(_08663_),
    .X(_08773_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15312_ (.A(_08773_),
    .X(_08774_));
 sky130_fd_sc_hd__a211o_1 _15313_ (.A1(_08231_),
    .A2(_08761_),
    .B1(_08772_),
    .C1(_08774_),
    .X(_08775_));
 sky130_fd_sc_hd__o22a_1 _15314_ (.A1(\irq_pending[1] ),
    .A2(_08542_),
    .B1(_08755_),
    .B2(_08775_),
    .X(_14583_));
 sky130_fd_sc_hd__mux2_1 _15315_ (.A0(\cpuregs[18][2] ),
    .A1(\cpuregs[19][2] ),
    .S(_08698_),
    .X(_08776_));
 sky130_fd_sc_hd__or2_1 _15316_ (.A(\cpuregs[16][2] ),
    .B(_08698_),
    .X(_08777_));
 sky130_fd_sc_hd__o211a_1 _15317_ (.A1(\cpuregs[17][2] ),
    .A2(_08700_),
    .B1(_08702_),
    .C1(_08777_),
    .X(_08778_));
 sky130_fd_sc_hd__a21oi_1 _15318_ (.A1(_08693_),
    .A2(_08776_),
    .B1(_08778_),
    .Y(_08779_));
 sky130_fd_sc_hd__mux2_1 _15319_ (.A0(\cpuregs[8][2] ),
    .A1(\cpuregs[9][2] ),
    .S(_08719_),
    .X(_08780_));
 sky130_fd_sc_hd__mux2_1 _15320_ (.A0(\cpuregs[10][2] ),
    .A1(\cpuregs[11][2] ),
    .S(_08719_),
    .X(_08781_));
 sky130_fd_sc_hd__mux2_1 _15321_ (.A0(_08780_),
    .A1(_08781_),
    .S(_08714_),
    .X(_08782_));
 sky130_fd_sc_hd__buf_2 _15322_ (.A(_08718_),
    .X(_08783_));
 sky130_fd_sc_hd__mux2_1 _15323_ (.A0(\cpuregs[12][2] ),
    .A1(\cpuregs[13][2] ),
    .S(_08783_),
    .X(_08784_));
 sky130_fd_sc_hd__mux2_1 _15324_ (.A0(\cpuregs[14][2] ),
    .A1(\cpuregs[15][2] ),
    .S(_08718_),
    .X(_08785_));
 sky130_fd_sc_hd__or2_1 _15325_ (.A(_08721_),
    .B(_08785_),
    .X(_08786_));
 sky130_fd_sc_hd__o211a_1 _15326_ (.A1(_08716_),
    .A2(_08784_),
    .B1(_08786_),
    .C1(_08724_),
    .X(_08787_));
 sky130_fd_sc_hd__a211o_1 _15327_ (.A1(_08708_),
    .A2(_08782_),
    .B1(_08787_),
    .C1(_08726_),
    .X(_08788_));
 sky130_fd_sc_hd__mux2_1 _15328_ (.A0(\cpuregs[2][2] ),
    .A1(\cpuregs[3][2] ),
    .S(_08710_),
    .X(_08789_));
 sky130_fd_sc_hd__or2_1 _15329_ (.A(_08732_),
    .B(_08789_),
    .X(_08790_));
 sky130_fd_sc_hd__mux2_1 _15330_ (.A0(\cpuregs[0][2] ),
    .A1(\cpuregs[1][2] ),
    .S(_08710_),
    .X(_08791_));
 sky130_fd_sc_hd__o21a_1 _15331_ (.A1(_08714_),
    .A2(_08791_),
    .B1(_08608_),
    .X(_08792_));
 sky130_fd_sc_hd__mux2_1 _15332_ (.A0(\cpuregs[6][2] ),
    .A1(\cpuregs[7][2] ),
    .S(_08560_),
    .X(_08793_));
 sky130_fd_sc_hd__mux2_1 _15333_ (.A0(\cpuregs[4][2] ),
    .A1(\cpuregs[5][2] ),
    .S(_08560_),
    .X(_08794_));
 sky130_fd_sc_hd__mux2_1 _15334_ (.A0(_08793_),
    .A1(_08794_),
    .S(_08569_),
    .X(_08795_));
 sky130_fd_sc_hd__a221o_1 _15335_ (.A1(_08790_),
    .A2(_08792_),
    .B1(_08795_),
    .B2(_08724_),
    .C1(_08740_),
    .X(_08796_));
 sky130_fd_sc_hd__a21oi_1 _15336_ (.A1(_08788_),
    .A2(_08796_),
    .B1(_08692_),
    .Y(_08797_));
 sky130_fd_sc_hd__a211o_4 _15337_ (.A1(_08692_),
    .A2(_08779_),
    .B1(_08797_),
    .C1(_08743_),
    .X(_08798_));
 sky130_fd_sc_hd__nor2_1 _15338_ (.A(_08690_),
    .B(_08798_),
    .Y(_08799_));
 sky130_fd_sc_hd__a221o_1 _15339_ (.A1(\irq_mask[2] ),
    .A2(_08639_),
    .B1(\timer[2] ),
    .B2(_08643_),
    .C1(_08647_),
    .X(_08800_));
 sky130_fd_sc_hd__buf_2 _15340_ (.A(instr_rdinstrh),
    .X(_08801_));
 sky130_fd_sc_hd__clkbuf_2 _15341_ (.A(_08801_),
    .X(_08802_));
 sky130_fd_sc_hd__clkbuf_2 _15342_ (.A(instr_rdinstr),
    .X(_08803_));
 sky130_fd_sc_hd__clkbuf_2 _15343_ (.A(instr_rdcycleh),
    .X(_08804_));
 sky130_fd_sc_hd__buf_2 _15344_ (.A(_08804_),
    .X(_08805_));
 sky130_fd_sc_hd__a22o_1 _15345_ (.A1(\count_instr[2] ),
    .A2(_08803_),
    .B1(_08805_),
    .B2(\count_cycle[34] ),
    .X(_08806_));
 sky130_fd_sc_hd__a21o_1 _15346_ (.A1(\count_instr[34] ),
    .A2(_08802_),
    .B1(_08806_),
    .X(_08807_));
 sky130_fd_sc_hd__a211o_1 _15347_ (.A1(\count_cycle[2] ),
    .A2(_08748_),
    .B1(_08807_),
    .C1(_08753_),
    .X(_08808_));
 sky130_fd_sc_hd__o211a_1 _15348_ (.A1(_08799_),
    .A2(_08800_),
    .B1(_08808_),
    .C1(_08181_),
    .X(_08809_));
 sky130_fd_sc_hd__clkbuf_2 _15349_ (.A(_08773_),
    .X(_08810_));
 sky130_fd_sc_hd__o211a_1 _15350_ (.A1(_08679_),
    .A2(net34),
    .B1(_08508_),
    .C1(_08191_),
    .X(_08811_));
 sky130_fd_sc_hd__o21a_1 _15351_ (.A1(net51),
    .A2(_08757_),
    .B1(_08811_),
    .X(_08812_));
 sky130_fd_sc_hd__a221o_1 _15352_ (.A1(net42),
    .A2(_08756_),
    .B1(_08678_),
    .B2(net55),
    .C1(_08812_),
    .X(_08813_));
 sky130_fd_sc_hd__mux2_2 _15353_ (.A0(\genblk1.pcpi_mul.rd[2] ),
    .A1(\genblk1.pcpi_mul.rd[34] ),
    .S(_08683_),
    .X(_08814_));
 sky130_fd_sc_hd__nand2_1 _15354_ (.A(\reg_pc[2] ),
    .B(\decoded_imm[2] ),
    .Y(_08815_));
 sky130_fd_sc_hd__or2_1 _15355_ (.A(\reg_pc[2] ),
    .B(\decoded_imm[2] ),
    .X(_08816_));
 sky130_fd_sc_hd__and2_1 _15356_ (.A(_08184_),
    .B(_08762_),
    .X(_08817_));
 sky130_fd_sc_hd__a31o_1 _15357_ (.A1(\reg_next_pc[0] ),
    .A2(\decoded_imm[0] ),
    .A3(_08764_),
    .B1(_08817_),
    .X(_08818_));
 sky130_fd_sc_hd__and3_1 _15358_ (.A(_08815_),
    .B(_08816_),
    .C(_08818_),
    .X(_08819_));
 sky130_fd_sc_hd__a21o_1 _15359_ (.A1(_08815_),
    .A2(_08816_),
    .B1(_08818_),
    .X(_08820_));
 sky130_fd_sc_hd__and3b_1 _15360_ (.A_N(_08819_),
    .B(_08820_),
    .C(_08311_),
    .X(_08821_));
 sky130_fd_sc_hd__a221o_1 _15361_ (.A1(_08671_),
    .A2(_08813_),
    .B1(_08814_),
    .B2(_08685_),
    .C1(_08821_),
    .X(_08822_));
 sky130_fd_sc_hd__or2_1 _15362_ (.A(_08810_),
    .B(_08822_),
    .X(_08823_));
 sky130_fd_sc_hd__o22a_1 _15363_ (.A1(\irq_pending[2] ),
    .A2(_08542_),
    .B1(_08809_),
    .B2(_08823_),
    .X(_14594_));
 sky130_fd_sc_hd__buf_2 _15364_ (.A(_08544_),
    .X(_08824_));
 sky130_fd_sc_hd__buf_2 _15365_ (.A(_08719_),
    .X(_08825_));
 sky130_fd_sc_hd__mux2_1 _15366_ (.A0(\cpuregs[16][3] ),
    .A1(\cpuregs[17][3] ),
    .S(_08825_),
    .X(_08826_));
 sky130_fd_sc_hd__clkbuf_2 _15367_ (.A(_08563_),
    .X(_08827_));
 sky130_fd_sc_hd__or2_1 _15368_ (.A(\cpuregs[18][3] ),
    .B(_08697_),
    .X(_08828_));
 sky130_fd_sc_hd__o211a_1 _15369_ (.A1(\cpuregs[19][3] ),
    .A2(_08827_),
    .B1(_08716_),
    .C1(_08828_),
    .X(_08829_));
 sky130_fd_sc_hd__a21oi_1 _15370_ (.A1(_08701_),
    .A2(_08826_),
    .B1(_08829_),
    .Y(_08830_));
 sky130_fd_sc_hd__buf_2 _15371_ (.A(_08580_),
    .X(_08831_));
 sky130_fd_sc_hd__buf_2 _15372_ (.A(_08556_),
    .X(_08832_));
 sky130_fd_sc_hd__clkbuf_4 _15373_ (.A(_08832_),
    .X(_08833_));
 sky130_fd_sc_hd__mux2_1 _15374_ (.A0(\cpuregs[8][3] ),
    .A1(\cpuregs[9][3] ),
    .S(_08833_),
    .X(_08834_));
 sky130_fd_sc_hd__clkbuf_4 _15375_ (.A(_08832_),
    .X(_08835_));
 sky130_fd_sc_hd__mux2_1 _15376_ (.A0(\cpuregs[10][3] ),
    .A1(\cpuregs[11][3] ),
    .S(_08835_),
    .X(_08836_));
 sky130_fd_sc_hd__clkbuf_4 _15377_ (.A(_08630_),
    .X(_08837_));
 sky130_fd_sc_hd__mux2_1 _15378_ (.A0(_08834_),
    .A1(_08836_),
    .S(_08837_),
    .X(_08838_));
 sky130_fd_sc_hd__buf_2 _15379_ (.A(_08588_),
    .X(_08839_));
 sky130_fd_sc_hd__buf_2 _15380_ (.A(_08571_),
    .X(_08840_));
 sky130_fd_sc_hd__mux2_1 _15381_ (.A0(\cpuregs[12][3] ),
    .A1(\cpuregs[13][3] ),
    .S(_08840_),
    .X(_08841_));
 sky130_fd_sc_hd__clkbuf_4 _15382_ (.A(_08557_),
    .X(_08842_));
 sky130_fd_sc_hd__mux2_1 _15383_ (.A0(\cpuregs[14][3] ),
    .A1(\cpuregs[15][3] ),
    .S(_08842_),
    .X(_08843_));
 sky130_fd_sc_hd__or2_1 _15384_ (.A(_08735_),
    .B(_08843_),
    .X(_08844_));
 sky130_fd_sc_hd__buf_2 _15385_ (.A(_08599_),
    .X(_08845_));
 sky130_fd_sc_hd__o211a_1 _15386_ (.A1(_08839_),
    .A2(_08841_),
    .B1(_08844_),
    .C1(_08845_),
    .X(_08846_));
 sky130_fd_sc_hd__buf_2 _15387_ (.A(_08604_),
    .X(_08847_));
 sky130_fd_sc_hd__a211o_1 _15388_ (.A1(_08831_),
    .A2(_08838_),
    .B1(_08846_),
    .C1(_08847_),
    .X(_08848_));
 sky130_fd_sc_hd__mux2_1 _15389_ (.A0(\cpuregs[2][3] ),
    .A1(\cpuregs[3][3] ),
    .S(_08559_),
    .X(_08849_));
 sky130_fd_sc_hd__or2_1 _15390_ (.A(_08731_),
    .B(_08849_),
    .X(_08850_));
 sky130_fd_sc_hd__clkbuf_4 _15391_ (.A(_08630_),
    .X(_08851_));
 sky130_fd_sc_hd__mux2_1 _15392_ (.A0(\cpuregs[0][3] ),
    .A1(\cpuregs[1][3] ),
    .S(_08835_),
    .X(_08852_));
 sky130_fd_sc_hd__o21a_1 _15393_ (.A1(_08851_),
    .A2(_08852_),
    .B1(_08706_),
    .X(_08853_));
 sky130_fd_sc_hd__buf_4 _15394_ (.A(_08694_),
    .X(_08854_));
 sky130_fd_sc_hd__mux2_1 _15395_ (.A0(\cpuregs[6][3] ),
    .A1(\cpuregs[7][3] ),
    .S(_08854_),
    .X(_08855_));
 sky130_fd_sc_hd__mux2_1 _15396_ (.A0(\cpuregs[4][3] ),
    .A1(\cpuregs[5][3] ),
    .S(_08854_),
    .X(_08856_));
 sky130_fd_sc_hd__clkbuf_4 _15397_ (.A(_08585_),
    .X(_08857_));
 sky130_fd_sc_hd__mux2_1 _15398_ (.A0(_08855_),
    .A1(_08856_),
    .S(_08857_),
    .X(_08858_));
 sky130_fd_sc_hd__buf_2 _15399_ (.A(_08598_),
    .X(_08859_));
 sky130_fd_sc_hd__clkbuf_4 _15400_ (.A(_08859_),
    .X(_08860_));
 sky130_fd_sc_hd__buf_2 _15401_ (.A(_08615_),
    .X(_08861_));
 sky130_fd_sc_hd__a221o_1 _15402_ (.A1(_08850_),
    .A2(_08853_),
    .B1(_08858_),
    .B2(_08860_),
    .C1(_08861_),
    .X(_08862_));
 sky130_fd_sc_hd__a21oi_2 _15403_ (.A1(_08848_),
    .A2(_08862_),
    .B1(_08691_),
    .Y(_08863_));
 sky130_fd_sc_hd__clkbuf_4 _15404_ (.A(_08632_),
    .X(_08864_));
 sky130_fd_sc_hd__a211o_4 _15405_ (.A1(_08824_),
    .A2(_08830_),
    .B1(_08863_),
    .C1(_08864_),
    .X(_08865_));
 sky130_fd_sc_hd__nor2_1 _15406_ (.A(_08690_),
    .B(_08865_),
    .Y(_08866_));
 sky130_fd_sc_hd__a221o_1 _15407_ (.A1(\irq_mask[3] ),
    .A2(_08639_),
    .B1(\timer[3] ),
    .B2(_08643_),
    .C1(_08647_),
    .X(_08867_));
 sky130_fd_sc_hd__a22o_1 _15408_ (.A1(\count_instr[3] ),
    .A2(_08803_),
    .B1(_08805_),
    .B2(\count_cycle[35] ),
    .X(_08868_));
 sky130_fd_sc_hd__a21o_1 _15409_ (.A1(\count_instr[35] ),
    .A2(_08802_),
    .B1(_08868_),
    .X(_08869_));
 sky130_fd_sc_hd__a211o_1 _15410_ (.A1(\count_cycle[3] ),
    .A2(_08748_),
    .B1(_08869_),
    .C1(_08753_),
    .X(_08870_));
 sky130_fd_sc_hd__o211a_1 _15411_ (.A1(_08866_),
    .A2(_08867_),
    .B1(_08870_),
    .C1(_08181_),
    .X(_08871_));
 sky130_fd_sc_hd__clkbuf_2 _15412_ (.A(_08312_),
    .X(_08872_));
 sky130_fd_sc_hd__clkbuf_2 _15413_ (.A(_08872_),
    .X(_08873_));
 sky130_fd_sc_hd__clkbuf_2 _15414_ (.A(\reg_pc[3] ),
    .X(_08874_));
 sky130_fd_sc_hd__nand2_1 _15415_ (.A(_08874_),
    .B(\decoded_imm[3] ),
    .Y(_08875_));
 sky130_fd_sc_hd__or2_1 _15416_ (.A(\reg_pc[3] ),
    .B(\decoded_imm[3] ),
    .X(_08876_));
 sky130_fd_sc_hd__nand2_1 _15417_ (.A(_08875_),
    .B(_08876_),
    .Y(_08877_));
 sky130_fd_sc_hd__a21bo_1 _15418_ (.A1(_08816_),
    .A2(_08818_),
    .B1_N(_08815_),
    .X(_08878_));
 sky130_fd_sc_hd__xnor2_1 _15419_ (.A(_08877_),
    .B(_08878_),
    .Y(_08879_));
 sky130_fd_sc_hd__clkbuf_2 _15420_ (.A(_08152_),
    .X(_08880_));
 sky130_fd_sc_hd__mux2_1 _15421_ (.A0(net35),
    .A1(net52),
    .S(_08679_),
    .X(_08881_));
 sky130_fd_sc_hd__and3_1 _15422_ (.A(_08325_),
    .B(_08509_),
    .C(_08881_),
    .X(_08882_));
 sky130_fd_sc_hd__a221o_1 _15423_ (.A1(net43),
    .A2(_08756_),
    .B1(net194),
    .B2(net58),
    .C1(_08882_),
    .X(_08883_));
 sky130_fd_sc_hd__buf_2 _15424_ (.A(_08768_),
    .X(_08884_));
 sky130_fd_sc_hd__mux2_2 _15425_ (.A0(\genblk1.pcpi_mul.rd[3] ),
    .A1(\genblk1.pcpi_mul.rd[35] ),
    .S(_08884_),
    .X(_08885_));
 sky130_fd_sc_hd__clkbuf_2 _15426_ (.A(_08287_),
    .X(_08886_));
 sky130_fd_sc_hd__a22o_1 _15427_ (.A1(_08880_),
    .A2(_08883_),
    .B1(_08885_),
    .B2(_08886_),
    .X(_08887_));
 sky130_fd_sc_hd__a211o_1 _15428_ (.A1(_08873_),
    .A2(_08879_),
    .B1(_08887_),
    .C1(_08774_),
    .X(_08888_));
 sky130_fd_sc_hd__o22a_1 _15429_ (.A1(\irq_pending[3] ),
    .A2(_08542_),
    .B1(_08871_),
    .B2(_08888_),
    .X(_14597_));
 sky130_fd_sc_hd__nand2_1 _15430_ (.A(\reg_pc[4] ),
    .B(\decoded_imm[4] ),
    .Y(_08889_));
 sky130_fd_sc_hd__or2_1 _15431_ (.A(\reg_pc[4] ),
    .B(\decoded_imm[4] ),
    .X(_08890_));
 sky130_fd_sc_hd__a21bo_1 _15432_ (.A1(_08876_),
    .A2(_08878_),
    .B1_N(_08875_),
    .X(_08891_));
 sky130_fd_sc_hd__and3_1 _15433_ (.A(_08889_),
    .B(_08890_),
    .C(_08891_),
    .X(_08892_));
 sky130_fd_sc_hd__a21o_1 _15434_ (.A1(_08889_),
    .A2(_08890_),
    .B1(_08891_),
    .X(_08893_));
 sky130_fd_sc_hd__clkbuf_2 _15435_ (.A(_08872_),
    .X(_08894_));
 sky130_fd_sc_hd__and3b_1 _15436_ (.A_N(_08892_),
    .B(_08893_),
    .C(_08894_),
    .X(_08895_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15437_ (.A(_08671_),
    .X(_08896_));
 sky130_fd_sc_hd__mux2_1 _15438_ (.A0(net36),
    .A1(net53),
    .S(_08758_),
    .X(_08897_));
 sky130_fd_sc_hd__and3_1 _15439_ (.A(_08326_),
    .B(_08509_),
    .C(_08897_),
    .X(_08898_));
 sky130_fd_sc_hd__a221o_1 _15440_ (.A1(net45),
    .A2(_08756_),
    .B1(net194),
    .B2(net59),
    .C1(_08898_),
    .X(_08899_));
 sky130_fd_sc_hd__buf_2 _15441_ (.A(_08683_),
    .X(_08900_));
 sky130_fd_sc_hd__mux2_4 _15442_ (.A0(\genblk1.pcpi_mul.rd[4] ),
    .A1(\genblk1.pcpi_mul.rd[36] ),
    .S(_08900_),
    .X(_08901_));
 sky130_fd_sc_hd__clkbuf_2 _15443_ (.A(_08288_),
    .X(_08902_));
 sky130_fd_sc_hd__clkbuf_4 _15444_ (.A(_08544_),
    .X(_08903_));
 sky130_fd_sc_hd__buf_2 _15445_ (.A(_08783_),
    .X(_08904_));
 sky130_fd_sc_hd__mux2_1 _15446_ (.A0(\cpuregs[16][4] ),
    .A1(\cpuregs[17][4] ),
    .S(_08904_),
    .X(_08905_));
 sky130_fd_sc_hd__or2_1 _15447_ (.A(\cpuregs[18][4] ),
    .B(_08629_),
    .X(_08906_));
 sky130_fd_sc_hd__o211a_1 _15448_ (.A1(\cpuregs[19][4] ),
    .A2(_08700_),
    .B1(_08552_),
    .C1(_08906_),
    .X(_08907_));
 sky130_fd_sc_hd__a21oi_1 _15449_ (.A1(_08702_),
    .A2(_08905_),
    .B1(_08907_),
    .Y(_08908_));
 sky130_fd_sc_hd__clkbuf_4 _15450_ (.A(_08595_),
    .X(_08909_));
 sky130_fd_sc_hd__mux2_1 _15451_ (.A0(\cpuregs[2][4] ),
    .A1(\cpuregs[3][4] ),
    .S(_08909_),
    .X(_08910_));
 sky130_fd_sc_hd__clkbuf_4 _15452_ (.A(_08594_),
    .X(_08911_));
 sky130_fd_sc_hd__clkbuf_4 _15453_ (.A(_08911_),
    .X(_08912_));
 sky130_fd_sc_hd__mux2_1 _15454_ (.A0(\cpuregs[0][4] ),
    .A1(\cpuregs[1][4] ),
    .S(_08912_),
    .X(_08913_));
 sky130_fd_sc_hd__mux2_1 _15455_ (.A0(_08910_),
    .A1(_08913_),
    .S(_08721_),
    .X(_08914_));
 sky130_fd_sc_hd__clkbuf_4 _15456_ (.A(_08550_),
    .X(_08915_));
 sky130_fd_sc_hd__mux2_1 _15457_ (.A0(\cpuregs[4][4] ),
    .A1(\cpuregs[5][4] ),
    .S(_08909_),
    .X(_08916_));
 sky130_fd_sc_hd__clkbuf_4 _15458_ (.A(_08567_),
    .X(_08917_));
 sky130_fd_sc_hd__buf_4 _15459_ (.A(_08594_),
    .X(_08918_));
 sky130_fd_sc_hd__mux2_1 _15460_ (.A0(\cpuregs[6][4] ),
    .A1(\cpuregs[7][4] ),
    .S(_08918_),
    .X(_08919_));
 sky130_fd_sc_hd__or2_1 _15461_ (.A(_08917_),
    .B(_08919_),
    .X(_08920_));
 sky130_fd_sc_hd__clkbuf_4 _15462_ (.A(_08599_),
    .X(_08921_));
 sky130_fd_sc_hd__o211a_1 _15463_ (.A1(_08915_),
    .A2(_08916_),
    .B1(_08920_),
    .C1(_08921_),
    .X(_08922_));
 sky130_fd_sc_hd__a211o_1 _15464_ (.A1(_08708_),
    .A2(_08914_),
    .B1(_08922_),
    .C1(_08740_),
    .X(_08923_));
 sky130_fd_sc_hd__mux2_1 _15465_ (.A0(\cpuregs[14][4] ),
    .A1(\cpuregs[15][4] ),
    .S(_08912_),
    .X(_08924_));
 sky130_fd_sc_hd__mux2_1 _15466_ (.A0(\cpuregs[12][4] ),
    .A1(\cpuregs[13][4] ),
    .S(_08912_),
    .X(_08925_));
 sky130_fd_sc_hd__mux2_1 _15467_ (.A0(_08924_),
    .A1(_08925_),
    .S(_08721_),
    .X(_08926_));
 sky130_fd_sc_hd__mux2_1 _15468_ (.A0(\cpuregs[8][4] ),
    .A1(\cpuregs[9][4] ),
    .S(_08909_),
    .X(_08927_));
 sky130_fd_sc_hd__mux2_1 _15469_ (.A0(\cpuregs[10][4] ),
    .A1(\cpuregs[11][4] ),
    .S(_08717_),
    .X(_08928_));
 sky130_fd_sc_hd__or2_1 _15470_ (.A(_08917_),
    .B(_08928_),
    .X(_08929_));
 sky130_fd_sc_hd__o211a_1 _15471_ (.A1(_08915_),
    .A2(_08927_),
    .B1(_08929_),
    .C1(_08707_),
    .X(_08930_));
 sky130_fd_sc_hd__a211o_1 _15472_ (.A1(_08724_),
    .A2(_08926_),
    .B1(_08930_),
    .C1(_08726_),
    .X(_08931_));
 sky130_fd_sc_hd__buf_4 _15473_ (.A(_08626_),
    .X(_08932_));
 sky130_fd_sc_hd__a21oi_1 _15474_ (.A1(_08923_),
    .A2(_08931_),
    .B1(_08932_),
    .Y(_08933_));
 sky130_fd_sc_hd__a211o_4 _15475_ (.A1(_08903_),
    .A2(_08908_),
    .B1(_08933_),
    .C1(_08743_),
    .X(_08934_));
 sky130_fd_sc_hd__nor2_1 _15476_ (.A(_08689_),
    .B(_08934_),
    .Y(_08935_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15477_ (.A(instr_maskirq),
    .X(_08936_));
 sky130_fd_sc_hd__clkbuf_2 _15478_ (.A(_08936_),
    .X(_08937_));
 sky130_fd_sc_hd__clkbuf_2 _15479_ (.A(_08640_),
    .X(_08938_));
 sky130_fd_sc_hd__clkbuf_2 _15480_ (.A(_08645_),
    .X(_08939_));
 sky130_fd_sc_hd__a221o_1 _15481_ (.A1(\irq_mask[4] ),
    .A2(_08937_),
    .B1(\timer[4] ),
    .B2(_08938_),
    .C1(_08939_),
    .X(_08940_));
 sky130_fd_sc_hd__clkbuf_2 _15482_ (.A(instr_rdinstr),
    .X(_08941_));
 sky130_fd_sc_hd__buf_2 _15483_ (.A(_08657_),
    .X(_08942_));
 sky130_fd_sc_hd__a22o_1 _15484_ (.A1(\count_instr[4] ),
    .A2(_08941_),
    .B1(_08942_),
    .B2(\count_instr[36] ),
    .X(_08943_));
 sky130_fd_sc_hd__a221o_1 _15485_ (.A1(_08652_),
    .A2(\count_cycle[36] ),
    .B1(_08747_),
    .B2(\count_cycle[4] ),
    .C1(_08943_),
    .X(_08944_));
 sky130_fd_sc_hd__clkbuf_4 _15486_ (.A(_08179_),
    .X(_08945_));
 sky130_fd_sc_hd__o221a_1 _15487_ (.A1(_08935_),
    .A2(_08940_),
    .B1(_08944_),
    .B2(_08752_),
    .C1(_08945_),
    .X(_08946_));
 sky130_fd_sc_hd__a221o_1 _15488_ (.A1(_08896_),
    .A2(_08899_),
    .B1(_08901_),
    .B2(_08902_),
    .C1(_08946_),
    .X(_08947_));
 sky130_fd_sc_hd__a211o_1 _15489_ (.A1(\irq_pending[4] ),
    .A2(_08774_),
    .B1(_08895_),
    .C1(_08947_),
    .X(_14598_));
 sky130_fd_sc_hd__buf_2 _15490_ (.A(_08714_),
    .X(_08948_));
 sky130_fd_sc_hd__mux2_1 _15491_ (.A0(\cpuregs[18][5] ),
    .A1(\cpuregs[19][5] ),
    .S(_08629_),
    .X(_08949_));
 sky130_fd_sc_hd__buf_2 _15492_ (.A(_08721_),
    .X(_08950_));
 sky130_fd_sc_hd__or2_1 _15493_ (.A(\cpuregs[16][5] ),
    .B(_08697_),
    .X(_08951_));
 sky130_fd_sc_hd__o211a_1 _15494_ (.A1(\cpuregs[17][5] ),
    .A2(_08827_),
    .B1(_08950_),
    .C1(_08951_),
    .X(_08952_));
 sky130_fd_sc_hd__a21oi_1 _15495_ (.A1(_08948_),
    .A2(_08949_),
    .B1(_08952_),
    .Y(_08953_));
 sky130_fd_sc_hd__clkbuf_4 _15496_ (.A(_08706_),
    .X(_08954_));
 sky130_fd_sc_hd__mux2_1 _15497_ (.A0(\cpuregs[2][5] ),
    .A1(\cpuregs[3][5] ),
    .S(_08709_),
    .X(_08955_));
 sky130_fd_sc_hd__mux2_1 _15498_ (.A0(\cpuregs[0][5] ),
    .A1(\cpuregs[1][5] ),
    .S(_08709_),
    .X(_08956_));
 sky130_fd_sc_hd__mux2_1 _15499_ (.A0(_08955_),
    .A1(_08956_),
    .S(_08857_),
    .X(_08957_));
 sky130_fd_sc_hd__mux2_1 _15500_ (.A0(\cpuregs[4][5] ),
    .A1(\cpuregs[5][5] ),
    .S(_08854_),
    .X(_08958_));
 sky130_fd_sc_hd__mux2_1 _15501_ (.A0(\cpuregs[6][5] ),
    .A1(\cpuregs[7][5] ),
    .S(_08558_),
    .X(_08959_));
 sky130_fd_sc_hd__or2_1 _15502_ (.A(_08730_),
    .B(_08959_),
    .X(_08960_));
 sky130_fd_sc_hd__o211a_1 _15503_ (.A1(_08837_),
    .A2(_08958_),
    .B1(_08960_),
    .C1(_08859_),
    .X(_08961_));
 sky130_fd_sc_hd__a211o_1 _15504_ (.A1(_08954_),
    .A2(_08957_),
    .B1(_08961_),
    .C1(_08861_),
    .X(_08962_));
 sky130_fd_sc_hd__buf_4 _15505_ (.A(_08594_),
    .X(_08963_));
 sky130_fd_sc_hd__mux2_1 _15506_ (.A0(\cpuregs[8][5] ),
    .A1(\cpuregs[9][5] ),
    .S(_08963_),
    .X(_08964_));
 sky130_fd_sc_hd__mux2_1 _15507_ (.A0(\cpuregs[10][5] ),
    .A1(\cpuregs[11][5] ),
    .S(_08963_),
    .X(_08965_));
 sky130_fd_sc_hd__mux2_1 _15508_ (.A0(_08964_),
    .A1(_08965_),
    .S(_08550_),
    .X(_08966_));
 sky130_fd_sc_hd__clkbuf_4 _15509_ (.A(_08630_),
    .X(_08967_));
 sky130_fd_sc_hd__mux2_1 _15510_ (.A0(\cpuregs[12][5] ),
    .A1(\cpuregs[13][5] ),
    .S(_08709_),
    .X(_08968_));
 sky130_fd_sc_hd__clkbuf_2 _15511_ (.A(_08592_),
    .X(_08969_));
 sky130_fd_sc_hd__clkbuf_2 _15512_ (.A(_08557_),
    .X(_08970_));
 sky130_fd_sc_hd__mux2_1 _15513_ (.A0(\cpuregs[14][5] ),
    .A1(\cpuregs[15][5] ),
    .S(_08970_),
    .X(_08971_));
 sky130_fd_sc_hd__or2_1 _15514_ (.A(_08969_),
    .B(_08971_),
    .X(_08972_));
 sky130_fd_sc_hd__buf_2 _15515_ (.A(_08598_),
    .X(_08973_));
 sky130_fd_sc_hd__o211a_1 _15516_ (.A1(_08967_),
    .A2(_08968_),
    .B1(_08972_),
    .C1(_08973_),
    .X(_08974_));
 sky130_fd_sc_hd__clkbuf_4 _15517_ (.A(_08603_),
    .X(_08975_));
 sky130_fd_sc_hd__a211o_1 _15518_ (.A1(_08954_),
    .A2(_08966_),
    .B1(_08974_),
    .C1(_08975_),
    .X(_08976_));
 sky130_fd_sc_hd__a21oi_2 _15519_ (.A1(_08962_),
    .A2(_08976_),
    .B1(_08691_),
    .Y(_08977_));
 sky130_fd_sc_hd__a211o_4 _15520_ (.A1(_08932_),
    .A2(_08953_),
    .B1(_08977_),
    .C1(_08864_),
    .X(_08978_));
 sky130_fd_sc_hd__nor2_1 _15521_ (.A(_08690_),
    .B(_08978_),
    .Y(_08979_));
 sky130_fd_sc_hd__a221o_1 _15522_ (.A1(\irq_mask[5] ),
    .A2(_08639_),
    .B1(\timer[5] ),
    .B2(_08643_),
    .C1(_08647_),
    .X(_08980_));
 sky130_fd_sc_hd__a22o_1 _15523_ (.A1(\count_instr[5] ),
    .A2(_08656_),
    .B1(_08805_),
    .B2(\count_cycle[37] ),
    .X(_08981_));
 sky130_fd_sc_hd__a21o_1 _15524_ (.A1(\count_instr[37] ),
    .A2(_08802_),
    .B1(_08981_),
    .X(_08982_));
 sky130_fd_sc_hd__a211o_1 _15525_ (.A1(\count_cycle[5] ),
    .A2(_08748_),
    .B1(_08982_),
    .C1(_08753_),
    .X(_08983_));
 sky130_fd_sc_hd__o211a_1 _15526_ (.A1(_08979_),
    .A2(_08980_),
    .B1(_08983_),
    .C1(_08181_),
    .X(_08984_));
 sky130_vsdinv _15527_ (.A(_08889_),
    .Y(_08985_));
 sky130_fd_sc_hd__or2_1 _15528_ (.A(_08985_),
    .B(_08892_),
    .X(_08986_));
 sky130_fd_sc_hd__nor2_1 _15529_ (.A(\reg_pc[5] ),
    .B(\decoded_imm[5] ),
    .Y(_08987_));
 sky130_fd_sc_hd__and2_1 _15530_ (.A(\reg_pc[5] ),
    .B(\decoded_imm[5] ),
    .X(_08988_));
 sky130_fd_sc_hd__or2_1 _15531_ (.A(_08987_),
    .B(_08988_),
    .X(_08989_));
 sky130_fd_sc_hd__xnor2_1 _15532_ (.A(_08986_),
    .B(_08989_),
    .Y(_08990_));
 sky130_fd_sc_hd__o211a_1 _15533_ (.A1(_08758_),
    .A2(net37),
    .B1(_08509_),
    .C1(_08325_),
    .X(_08991_));
 sky130_fd_sc_hd__o21a_1 _15534_ (.A1(_08757_),
    .A2(net54),
    .B1(_08991_),
    .X(_08992_));
 sky130_fd_sc_hd__a221o_1 _15535_ (.A1(net46),
    .A2(_08756_),
    .B1(net194),
    .B2(net60),
    .C1(_08992_),
    .X(_08993_));
 sky130_fd_sc_hd__mux2_2 _15536_ (.A0(\genblk1.pcpi_mul.rd[5] ),
    .A1(\genblk1.pcpi_mul.rd[37] ),
    .S(_08884_),
    .X(_08994_));
 sky130_fd_sc_hd__a22o_1 _15537_ (.A1(_08880_),
    .A2(_08993_),
    .B1(_08994_),
    .B2(_08886_),
    .X(_08995_));
 sky130_fd_sc_hd__a211o_1 _15538_ (.A1(_08894_),
    .A2(_08990_),
    .B1(_08995_),
    .C1(_08810_),
    .X(_08996_));
 sky130_fd_sc_hd__o22a_1 _15539_ (.A1(\irq_pending[5] ),
    .A2(_08542_),
    .B1(_08984_),
    .B2(_08996_),
    .X(_14599_));
 sky130_fd_sc_hd__clkbuf_2 _15540_ (.A(\reg_pc[6] ),
    .X(_08997_));
 sky130_fd_sc_hd__nand2_1 _15541_ (.A(_08997_),
    .B(\decoded_imm[6] ),
    .Y(_08998_));
 sky130_fd_sc_hd__or2_1 _15542_ (.A(\reg_pc[6] ),
    .B(\decoded_imm[6] ),
    .X(_08999_));
 sky130_fd_sc_hd__nand2_1 _15543_ (.A(_08998_),
    .B(_08999_),
    .Y(_09000_));
 sky130_fd_sc_hd__a211oi_1 _15544_ (.A1(_08890_),
    .A2(_08891_),
    .B1(_08988_),
    .C1(_08985_),
    .Y(_09001_));
 sky130_fd_sc_hd__nor2_1 _15545_ (.A(_08987_),
    .B(_09001_),
    .Y(_09002_));
 sky130_fd_sc_hd__xnor2_1 _15546_ (.A(_09000_),
    .B(_09002_),
    .Y(_09003_));
 sky130_fd_sc_hd__o211a_1 _15547_ (.A1(_08679_),
    .A2(net38),
    .B1(_08508_),
    .C1(_08191_),
    .X(_09004_));
 sky130_fd_sc_hd__o21a_1 _15548_ (.A1(_08757_),
    .A2(net56),
    .B1(_09004_),
    .X(_09005_));
 sky130_fd_sc_hd__a221o_1 _15549_ (.A1(net47),
    .A2(_08756_),
    .B1(_08678_),
    .B2(net61),
    .C1(_09005_),
    .X(_09006_));
 sky130_fd_sc_hd__mux2_2 _15550_ (.A0(\genblk1.pcpi_mul.rd[6] ),
    .A1(\genblk1.pcpi_mul.rd[38] ),
    .S(_08769_),
    .X(_09007_));
 sky130_fd_sc_hd__a22o_1 _15551_ (.A1(_08880_),
    .A2(_09006_),
    .B1(_09007_),
    .B2(_08288_),
    .X(_09008_));
 sky130_fd_sc_hd__clkbuf_2 _15552_ (.A(_08689_),
    .X(_09009_));
 sky130_fd_sc_hd__mux2_1 _15553_ (.A0(\cpuregs[16][6] ),
    .A1(\cpuregs[17][6] ),
    .S(_08698_),
    .X(_09010_));
 sky130_fd_sc_hd__or2_1 _15554_ (.A(\cpuregs[18][6] ),
    .B(_08904_),
    .X(_09011_));
 sky130_fd_sc_hd__o211a_1 _15555_ (.A1(\cpuregs[19][6] ),
    .A2(_08700_),
    .B1(_08948_),
    .C1(_09011_),
    .X(_09012_));
 sky130_fd_sc_hd__a21oi_1 _15556_ (.A1(_08702_),
    .A2(_09010_),
    .B1(_09012_),
    .Y(_09013_));
 sky130_fd_sc_hd__mux2_1 _15557_ (.A0(\cpuregs[8][6] ),
    .A1(\cpuregs[9][6] ),
    .S(_08573_),
    .X(_09014_));
 sky130_fd_sc_hd__mux2_1 _15558_ (.A0(\cpuregs[10][6] ),
    .A1(\cpuregs[11][6] ),
    .S(_08573_),
    .X(_09015_));
 sky130_fd_sc_hd__mux2_1 _15559_ (.A0(_09014_),
    .A1(_09015_),
    .S(_08915_),
    .X(_09016_));
 sky130_fd_sc_hd__mux2_1 _15560_ (.A0(\cpuregs[12][6] ),
    .A1(\cpuregs[13][6] ),
    .S(_08573_),
    .X(_09017_));
 sky130_fd_sc_hd__clkbuf_4 _15561_ (.A(_08969_),
    .X(_09018_));
 sky130_fd_sc_hd__mux2_1 _15562_ (.A0(\cpuregs[14][6] ),
    .A1(\cpuregs[15][6] ),
    .S(_08854_),
    .X(_09019_));
 sky130_fd_sc_hd__or2_1 _15563_ (.A(_09018_),
    .B(_09019_),
    .X(_09020_));
 sky130_fd_sc_hd__o211a_1 _15564_ (.A1(_08714_),
    .A2(_09017_),
    .B1(_09020_),
    .C1(_08921_),
    .X(_09021_));
 sky130_fd_sc_hd__a211o_1 _15565_ (.A1(_08708_),
    .A2(_09016_),
    .B1(_09021_),
    .C1(_08726_),
    .X(_09022_));
 sky130_fd_sc_hd__mux2_1 _15566_ (.A0(\cpuregs[2][6] ),
    .A1(\cpuregs[3][6] ),
    .S(_08696_),
    .X(_09023_));
 sky130_fd_sc_hd__or2_1 _15567_ (.A(_08569_),
    .B(_09023_),
    .X(_09024_));
 sky130_fd_sc_hd__mux2_1 _15568_ (.A0(\cpuregs[0][6] ),
    .A1(\cpuregs[1][6] ),
    .S(_08696_),
    .X(_09025_));
 sky130_fd_sc_hd__clkbuf_4 _15569_ (.A(_08706_),
    .X(_09026_));
 sky130_fd_sc_hd__o21a_1 _15570_ (.A1(_08714_),
    .A2(_09025_),
    .B1(_09026_),
    .X(_09027_));
 sky130_fd_sc_hd__mux2_1 _15571_ (.A0(\cpuregs[6][6] ),
    .A1(\cpuregs[7][6] ),
    .S(_08696_),
    .X(_09028_));
 sky130_fd_sc_hd__mux2_1 _15572_ (.A0(\cpuregs[4][6] ),
    .A1(\cpuregs[5][6] ),
    .S(_08696_),
    .X(_09029_));
 sky130_fd_sc_hd__mux2_1 _15573_ (.A0(_09028_),
    .A1(_09029_),
    .S(_08569_),
    .X(_09030_));
 sky130_fd_sc_hd__a221o_1 _15574_ (.A1(_09024_),
    .A2(_09027_),
    .B1(_09030_),
    .B2(_08724_),
    .C1(_08740_),
    .X(_09031_));
 sky130_fd_sc_hd__a21oi_1 _15575_ (.A1(_09022_),
    .A2(_09031_),
    .B1(_08903_),
    .Y(_09032_));
 sky130_fd_sc_hd__a211o_4 _15576_ (.A1(_08692_),
    .A2(_09013_),
    .B1(_09032_),
    .C1(_08743_),
    .X(_09033_));
 sky130_fd_sc_hd__nor2_1 _15577_ (.A(_09009_),
    .B(_09033_),
    .Y(_09034_));
 sky130_fd_sc_hd__clkbuf_2 _15578_ (.A(_08645_),
    .X(_09035_));
 sky130_fd_sc_hd__a221o_1 _15579_ (.A1(\irq_mask[6] ),
    .A2(_08638_),
    .B1(\timer[6] ),
    .B2(_08642_),
    .C1(_09035_),
    .X(_09036_));
 sky130_fd_sc_hd__clkbuf_2 _15580_ (.A(_08653_),
    .X(_09037_));
 sky130_fd_sc_hd__a22o_1 _15581_ (.A1(\count_instr[6] ),
    .A2(_08941_),
    .B1(_08804_),
    .B2(\count_cycle[38] ),
    .X(_09038_));
 sky130_fd_sc_hd__a21o_1 _15582_ (.A1(\count_instr[38] ),
    .A2(_08658_),
    .B1(_09038_),
    .X(_09039_));
 sky130_fd_sc_hd__a211o_1 _15583_ (.A1(\count_cycle[6] ),
    .A2(_09037_),
    .B1(_09039_),
    .C1(_08752_),
    .X(_09040_));
 sky130_fd_sc_hd__o211a_1 _15584_ (.A1(_09034_),
    .A2(_09036_),
    .B1(_09040_),
    .C1(_08293_),
    .X(_09041_));
 sky130_fd_sc_hd__a2111o_1 _15585_ (.A1(_08894_),
    .A2(_09003_),
    .B1(_09008_),
    .C1(_08810_),
    .D1(_09041_),
    .X(_09042_));
 sky130_fd_sc_hd__o21a_1 _15586_ (.A1(\irq_pending[6] ),
    .A2(_08542_),
    .B1(_09042_),
    .X(_14600_));
 sky130_fd_sc_hd__and2_1 _15587_ (.A(\reg_pc[7] ),
    .B(\decoded_imm[7] ),
    .X(_09043_));
 sky130_fd_sc_hd__nor2_1 _15588_ (.A(\reg_pc[7] ),
    .B(\decoded_imm[7] ),
    .Y(_09044_));
 sky130_fd_sc_hd__or2_1 _15589_ (.A(_09043_),
    .B(_09044_),
    .X(_09045_));
 sky130_fd_sc_hd__o31ai_1 _15590_ (.A1(_08987_),
    .A2(_09000_),
    .A3(_09001_),
    .B1(_08998_),
    .Y(_09046_));
 sky130_fd_sc_hd__xnor2_1 _15591_ (.A(_09045_),
    .B(_09046_),
    .Y(_09047_));
 sky130_fd_sc_hd__clkbuf_2 _15592_ (.A(_08671_),
    .X(_09048_));
 sky130_fd_sc_hd__or2_1 _15593_ (.A(_08672_),
    .B(net57),
    .X(_09049_));
 sky130_fd_sc_hd__o2111a_1 _15594_ (.A1(_08193_),
    .A2(net39),
    .B1(_09049_),
    .C1(_08508_),
    .D1(_08191_),
    .X(_09050_));
 sky130_fd_sc_hd__a221o_1 _15595_ (.A1(net48),
    .A2(_08675_),
    .B1(_08678_),
    .B2(net62),
    .C1(_09050_),
    .X(_09051_));
 sky130_fd_sc_hd__buf_2 _15596_ (.A(_08768_),
    .X(_09052_));
 sky130_fd_sc_hd__mux2_4 _15597_ (.A0(\genblk1.pcpi_mul.rd[7] ),
    .A1(\genblk1.pcpi_mul.rd[39] ),
    .S(_09052_),
    .X(_09053_));
 sky130_fd_sc_hd__mux2_1 _15598_ (.A0(\cpuregs[18][7] ),
    .A1(\cpuregs[19][7] ),
    .S(_08825_),
    .X(_09054_));
 sky130_fd_sc_hd__buf_2 _15599_ (.A(_08564_),
    .X(_09055_));
 sky130_fd_sc_hd__clkbuf_2 _15600_ (.A(_08573_),
    .X(_09056_));
 sky130_fd_sc_hd__or2_1 _15601_ (.A(\cpuregs[16][7] ),
    .B(_09056_),
    .X(_09057_));
 sky130_fd_sc_hd__o211a_1 _15602_ (.A1(\cpuregs[17][7] ),
    .A2(_09055_),
    .B1(_08950_),
    .C1(_09057_),
    .X(_09058_));
 sky130_fd_sc_hd__a21oi_1 _15603_ (.A1(_08553_),
    .A2(_09054_),
    .B1(_09058_),
    .Y(_09059_));
 sky130_fd_sc_hd__buf_4 _15604_ (.A(_08832_),
    .X(_09060_));
 sky130_fd_sc_hd__mux2_1 _15605_ (.A0(\cpuregs[10][7] ),
    .A1(\cpuregs[11][7] ),
    .S(_09060_),
    .X(_09061_));
 sky130_fd_sc_hd__buf_4 _15606_ (.A(_08832_),
    .X(_09062_));
 sky130_fd_sc_hd__mux2_1 _15607_ (.A0(\cpuregs[8][7] ),
    .A1(\cpuregs[9][7] ),
    .S(_09062_),
    .X(_09063_));
 sky130_fd_sc_hd__mux2_1 _15608_ (.A0(_09061_),
    .A1(_09063_),
    .S(_08613_),
    .X(_09064_));
 sky130_fd_sc_hd__buf_2 _15609_ (.A(_08588_),
    .X(_09065_));
 sky130_fd_sc_hd__clkbuf_4 _15610_ (.A(_08558_),
    .X(_09066_));
 sky130_fd_sc_hd__mux2_1 _15611_ (.A0(\cpuregs[12][7] ),
    .A1(\cpuregs[13][7] ),
    .S(_09066_),
    .X(_09067_));
 sky130_fd_sc_hd__clkbuf_2 _15612_ (.A(_08592_),
    .X(_09068_));
 sky130_fd_sc_hd__clkbuf_4 _15613_ (.A(_08557_),
    .X(_09069_));
 sky130_fd_sc_hd__mux2_1 _15614_ (.A0(\cpuregs[14][7] ),
    .A1(\cpuregs[15][7] ),
    .S(_09069_),
    .X(_09070_));
 sky130_fd_sc_hd__or2_1 _15615_ (.A(_09068_),
    .B(_09070_),
    .X(_09071_));
 sky130_fd_sc_hd__o211a_1 _15616_ (.A1(_09065_),
    .A2(_09067_),
    .B1(_09071_),
    .C1(_08845_),
    .X(_09072_));
 sky130_fd_sc_hd__buf_2 _15617_ (.A(_08604_),
    .X(_09073_));
 sky130_fd_sc_hd__a211o_1 _15618_ (.A1(_08831_),
    .A2(_09064_),
    .B1(_09072_),
    .C1(_09073_),
    .X(_09074_));
 sky130_fd_sc_hd__buf_2 _15619_ (.A(_08607_),
    .X(_09075_));
 sky130_fd_sc_hd__clkbuf_4 _15620_ (.A(_08609_),
    .X(_09076_));
 sky130_fd_sc_hd__mux2_1 _15621_ (.A0(\cpuregs[2][7] ),
    .A1(\cpuregs[3][7] ),
    .S(_09076_),
    .X(_09077_));
 sky130_fd_sc_hd__clkbuf_4 _15622_ (.A(_08609_),
    .X(_09078_));
 sky130_fd_sc_hd__mux2_1 _15623_ (.A0(\cpuregs[0][7] ),
    .A1(\cpuregs[1][7] ),
    .S(_09078_),
    .X(_09079_));
 sky130_fd_sc_hd__clkbuf_4 _15624_ (.A(_08567_),
    .X(_09080_));
 sky130_fd_sc_hd__mux2_1 _15625_ (.A0(_09077_),
    .A1(_09079_),
    .S(_09080_),
    .X(_09081_));
 sky130_fd_sc_hd__buf_2 _15626_ (.A(_08630_),
    .X(_09082_));
 sky130_fd_sc_hd__clkbuf_4 _15627_ (.A(_08970_),
    .X(_09083_));
 sky130_fd_sc_hd__mux2_1 _15628_ (.A0(\cpuregs[4][7] ),
    .A1(\cpuregs[5][7] ),
    .S(_09083_),
    .X(_09084_));
 sky130_fd_sc_hd__mux2_1 _15629_ (.A0(\cpuregs[6][7] ),
    .A1(\cpuregs[7][7] ),
    .S(_08911_),
    .X(_09085_));
 sky130_fd_sc_hd__or2_1 _15630_ (.A(_08730_),
    .B(_09085_),
    .X(_09086_));
 sky130_fd_sc_hd__buf_2 _15631_ (.A(_08598_),
    .X(_09087_));
 sky130_fd_sc_hd__o211a_1 _15632_ (.A1(_09082_),
    .A2(_09084_),
    .B1(_09086_),
    .C1(_09087_),
    .X(_09088_));
 sky130_fd_sc_hd__a211o_1 _15633_ (.A1(_09075_),
    .A2(_09081_),
    .B1(_09088_),
    .C1(_08617_),
    .X(_09089_));
 sky130_fd_sc_hd__buf_4 _15634_ (.A(_08543_),
    .X(_09090_));
 sky130_fd_sc_hd__a21oi_2 _15635_ (.A1(_09074_),
    .A2(_09089_),
    .B1(_09090_),
    .Y(_09091_));
 sky130_fd_sc_hd__clkbuf_4 _15636_ (.A(_08633_),
    .X(_09092_));
 sky130_fd_sc_hd__a211o_4 _15637_ (.A1(_08824_),
    .A2(_09059_),
    .B1(_09091_),
    .C1(_09092_),
    .X(_09093_));
 sky130_fd_sc_hd__nor2_1 _15638_ (.A(_08689_),
    .B(_09093_),
    .Y(_09094_));
 sky130_fd_sc_hd__clkbuf_2 _15639_ (.A(_08645_),
    .X(_09095_));
 sky130_fd_sc_hd__a221o_1 _15640_ (.A1(\irq_mask[7] ),
    .A2(_08937_),
    .B1(\timer[7] ),
    .B2(_08938_),
    .C1(_09095_),
    .X(_09096_));
 sky130_fd_sc_hd__a22o_1 _15641_ (.A1(\count_instr[39] ),
    .A2(_08657_),
    .B1(_08651_),
    .B2(\count_cycle[39] ),
    .X(_09097_));
 sky130_fd_sc_hd__a221o_1 _15642_ (.A1(\count_instr[7] ),
    .A2(_08803_),
    .B1(\count_cycle[7] ),
    .B2(_08747_),
    .C1(_09097_),
    .X(_09098_));
 sky130_fd_sc_hd__o221a_1 _15643_ (.A1(_09094_),
    .A2(_09096_),
    .B1(_09098_),
    .B2(_08752_),
    .C1(_08945_),
    .X(_09099_));
 sky130_fd_sc_hd__a221o_1 _15644_ (.A1(_09048_),
    .A2(_09051_),
    .B1(_09053_),
    .B2(_08517_),
    .C1(_09099_),
    .X(_09100_));
 sky130_fd_sc_hd__a221o_1 _15645_ (.A1(\irq_pending[7] ),
    .A2(_08774_),
    .B1(_09047_),
    .B2(_08873_),
    .C1(_09100_),
    .X(_14601_));
 sky130_fd_sc_hd__clkbuf_2 _15646_ (.A(_08873_),
    .X(_09101_));
 sky130_fd_sc_hd__or2_1 _15647_ (.A(\reg_pc[8] ),
    .B(\decoded_imm[8] ),
    .X(_09102_));
 sky130_fd_sc_hd__nand2_1 _15648_ (.A(\reg_pc[8] ),
    .B(\decoded_imm[8] ),
    .Y(_09103_));
 sky130_fd_sc_hd__and2b_1 _15649_ (.A_N(_09045_),
    .B(_09046_),
    .X(_09104_));
 sky130_fd_sc_hd__a211o_1 _15650_ (.A1(_09102_),
    .A2(_09103_),
    .B1(_09043_),
    .C1(_09104_),
    .X(_09105_));
 sky130_fd_sc_hd__o211ai_1 _15651_ (.A1(_09043_),
    .A2(_09104_),
    .B1(_09102_),
    .C1(_09103_),
    .Y(_09106_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15652_ (.A(_08540_),
    .X(_09107_));
 sky130_fd_sc_hd__clkbuf_4 _15653_ (.A(_08626_),
    .X(_09108_));
 sky130_fd_sc_hd__clkbuf_2 _15654_ (.A(_08570_),
    .X(_09109_));
 sky130_fd_sc_hd__clkbuf_4 _15655_ (.A(_08560_),
    .X(_09110_));
 sky130_fd_sc_hd__mux2_1 _15656_ (.A0(\cpuregs[16][8] ),
    .A1(\cpuregs[17][8] ),
    .S(_09110_),
    .X(_09111_));
 sky130_fd_sc_hd__buf_2 _15657_ (.A(_08564_),
    .X(_09112_));
 sky130_fd_sc_hd__clkbuf_2 _15658_ (.A(_08551_),
    .X(_09113_));
 sky130_fd_sc_hd__or2_1 _15659_ (.A(\cpuregs[18][8] ),
    .B(_09056_),
    .X(_09114_));
 sky130_fd_sc_hd__o211a_1 _15660_ (.A1(\cpuregs[19][8] ),
    .A2(_09112_),
    .B1(_09113_),
    .C1(_09114_),
    .X(_09115_));
 sky130_fd_sc_hd__a21oi_1 _15661_ (.A1(_09109_),
    .A2(_09111_),
    .B1(_09115_),
    .Y(_09116_));
 sky130_fd_sc_hd__buf_2 _15662_ (.A(_08580_),
    .X(_09117_));
 sky130_fd_sc_hd__buf_4 _15663_ (.A(_08970_),
    .X(_09118_));
 sky130_fd_sc_hd__mux2_1 _15664_ (.A0(\cpuregs[2][8] ),
    .A1(\cpuregs[3][8] ),
    .S(_09118_),
    .X(_09119_));
 sky130_fd_sc_hd__mux2_1 _15665_ (.A0(\cpuregs[0][8] ),
    .A1(\cpuregs[1][8] ),
    .S(_09060_),
    .X(_09120_));
 sky130_fd_sc_hd__clkbuf_4 _15666_ (.A(_08585_),
    .X(_09121_));
 sky130_fd_sc_hd__mux2_1 _15667_ (.A0(_09119_),
    .A1(_09120_),
    .S(_09121_),
    .X(_09122_));
 sky130_fd_sc_hd__buf_2 _15668_ (.A(_08588_),
    .X(_09123_));
 sky130_fd_sc_hd__clkbuf_4 _15669_ (.A(_08558_),
    .X(_09124_));
 sky130_fd_sc_hd__mux2_1 _15670_ (.A0(\cpuregs[4][8] ),
    .A1(\cpuregs[5][8] ),
    .S(_09124_),
    .X(_09125_));
 sky130_fd_sc_hd__clkbuf_2 _15671_ (.A(_08567_),
    .X(_09126_));
 sky130_fd_sc_hd__buf_4 _15672_ (.A(_08557_),
    .X(_09127_));
 sky130_fd_sc_hd__mux2_1 _15673_ (.A0(\cpuregs[6][8] ),
    .A1(\cpuregs[7][8] ),
    .S(_09127_),
    .X(_09128_));
 sky130_fd_sc_hd__or2_1 _15674_ (.A(_09126_),
    .B(_09128_),
    .X(_09129_));
 sky130_fd_sc_hd__buf_2 _15675_ (.A(_08599_),
    .X(_09130_));
 sky130_fd_sc_hd__o211a_1 _15676_ (.A1(_09123_),
    .A2(_09125_),
    .B1(_09129_),
    .C1(_09130_),
    .X(_09131_));
 sky130_fd_sc_hd__clkbuf_4 _15677_ (.A(_08616_),
    .X(_09132_));
 sky130_fd_sc_hd__a211o_1 _15678_ (.A1(_09117_),
    .A2(_09122_),
    .B1(_09131_),
    .C1(_09132_),
    .X(_09133_));
 sky130_fd_sc_hd__clkbuf_4 _15679_ (.A(_08609_),
    .X(_09134_));
 sky130_fd_sc_hd__mux2_1 _15680_ (.A0(\cpuregs[14][8] ),
    .A1(\cpuregs[15][8] ),
    .S(_09134_),
    .X(_09135_));
 sky130_fd_sc_hd__clkbuf_4 _15681_ (.A(_08609_),
    .X(_09136_));
 sky130_fd_sc_hd__mux2_1 _15682_ (.A0(\cpuregs[12][8] ),
    .A1(\cpuregs[13][8] ),
    .S(_09136_),
    .X(_09137_));
 sky130_fd_sc_hd__mux2_1 _15683_ (.A0(_09135_),
    .A1(_09137_),
    .S(_09080_),
    .X(_09138_));
 sky130_fd_sc_hd__buf_2 _15684_ (.A(_08588_),
    .X(_09139_));
 sky130_fd_sc_hd__clkbuf_4 _15685_ (.A(_08970_),
    .X(_09140_));
 sky130_fd_sc_hd__mux2_1 _15686_ (.A0(\cpuregs[8][8] ),
    .A1(\cpuregs[9][8] ),
    .S(_09140_),
    .X(_09141_));
 sky130_fd_sc_hd__clkbuf_2 _15687_ (.A(_08592_),
    .X(_09142_));
 sky130_fd_sc_hd__clkbuf_4 _15688_ (.A(_08556_),
    .X(_09143_));
 sky130_fd_sc_hd__mux2_1 _15689_ (.A0(\cpuregs[10][8] ),
    .A1(\cpuregs[11][8] ),
    .S(_09143_),
    .X(_09144_));
 sky130_fd_sc_hd__or2_1 _15690_ (.A(_09142_),
    .B(_09144_),
    .X(_09145_));
 sky130_fd_sc_hd__o211a_1 _15691_ (.A1(_09139_),
    .A2(_09141_),
    .B1(_09145_),
    .C1(_08607_),
    .X(_09146_));
 sky130_fd_sc_hd__a211o_1 _15692_ (.A1(_08860_),
    .A2(_09138_),
    .B1(_09146_),
    .C1(_08847_),
    .X(_09147_));
 sky130_fd_sc_hd__clkbuf_4 _15693_ (.A(_08626_),
    .X(_09148_));
 sky130_fd_sc_hd__a21oi_2 _15694_ (.A1(_09133_),
    .A2(_09147_),
    .B1(_09148_),
    .Y(_09149_));
 sky130_fd_sc_hd__clkbuf_4 _15695_ (.A(_08633_),
    .X(_09150_));
 sky130_fd_sc_hd__a211o_4 _15696_ (.A1(_09108_),
    .A2(_09116_),
    .B1(_09149_),
    .C1(_09150_),
    .X(_09151_));
 sky130_fd_sc_hd__nor2_1 _15697_ (.A(_09009_),
    .B(_09151_),
    .Y(_09152_));
 sky130_fd_sc_hd__a221o_1 _15698_ (.A1(\irq_mask[8] ),
    .A2(_08638_),
    .B1(\timer[8] ),
    .B2(_08642_),
    .C1(_08647_),
    .X(_09153_));
 sky130_fd_sc_hd__a22o_1 _15699_ (.A1(\count_instr[8] ),
    .A2(_08941_),
    .B1(_08651_),
    .B2(\count_cycle[40] ),
    .X(_09154_));
 sky130_fd_sc_hd__a21o_1 _15700_ (.A1(\count_instr[40] ),
    .A2(_08658_),
    .B1(_09154_),
    .X(_09155_));
 sky130_fd_sc_hd__a211o_1 _15701_ (.A1(\count_cycle[8] ),
    .A2(_09037_),
    .B1(_09155_),
    .C1(_08752_),
    .X(_09156_));
 sky130_fd_sc_hd__o211a_1 _15702_ (.A1(_09152_),
    .A2(_09153_),
    .B1(_09156_),
    .C1(_08180_),
    .X(_09157_));
 sky130_fd_sc_hd__mux2_4 _15703_ (.A0(\genblk1.pcpi_mul.rd[8] ),
    .A1(\genblk1.pcpi_mul.rd[40] ),
    .S(_09052_),
    .X(_09158_));
 sky130_fd_sc_hd__and2_1 _15704_ (.A(latched_is_lb),
    .B(_09051_),
    .X(_09159_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15705_ (.A(_09159_),
    .X(_09160_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15706_ (.A(_08674_),
    .X(_09161_));
 sky130_vsdinv _15707_ (.A(latched_is_lb),
    .Y(_09162_));
 sky130_fd_sc_hd__o21a_1 _15708_ (.A1(_09162_),
    .A2(latched_is_lh),
    .B1(_08677_),
    .X(_09163_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15709_ (.A(_09163_),
    .X(_09164_));
 sky130_fd_sc_hd__o221a_1 _15710_ (.A1(net63),
    .A2(_09161_),
    .B1(_08676_),
    .B2(net49),
    .C1(_09164_),
    .X(_09165_));
 sky130_fd_sc_hd__o21a_1 _15711_ (.A1(_09160_),
    .A2(_09165_),
    .B1(_08152_),
    .X(_09166_));
 sky130_fd_sc_hd__a211o_1 _15712_ (.A1(_08517_),
    .A2(_09158_),
    .B1(_09166_),
    .C1(_08773_),
    .X(_09167_));
 sky130_fd_sc_hd__o22a_1 _15713_ (.A1(\irq_pending[8] ),
    .A2(_09107_),
    .B1(_09157_),
    .B2(_09167_),
    .X(_09168_));
 sky130_fd_sc_hd__a31o_1 _15714_ (.A1(_09101_),
    .A2(_09105_),
    .A3(_09106_),
    .B1(_09168_),
    .X(_14602_));
 sky130_fd_sc_hd__or2_1 _15715_ (.A(\reg_pc[9] ),
    .B(\decoded_imm[9] ),
    .X(_09169_));
 sky130_fd_sc_hd__clkbuf_2 _15716_ (.A(\reg_pc[9] ),
    .X(_09170_));
 sky130_fd_sc_hd__nand2_1 _15717_ (.A(_09170_),
    .B(\decoded_imm[9] ),
    .Y(_09171_));
 sky130_fd_sc_hd__nand2_1 _15718_ (.A(_09169_),
    .B(_09171_),
    .Y(_09172_));
 sky130_fd_sc_hd__nand3_1 _15719_ (.A(_09103_),
    .B(_09106_),
    .C(_09172_),
    .Y(_09173_));
 sky130_vsdinv _15720_ (.A(_09172_),
    .Y(_09174_));
 sky130_fd_sc_hd__o2111ai_2 _15721_ (.A1(_09043_),
    .A2(_09104_),
    .B1(_09102_),
    .C1(_09103_),
    .D1(_09174_),
    .Y(_09175_));
 sky130_fd_sc_hd__or2_1 _15722_ (.A(_09103_),
    .B(_09172_),
    .X(_09176_));
 sky130_fd_sc_hd__and4_1 _15723_ (.A(_08872_),
    .B(_09173_),
    .C(_09175_),
    .D(_09176_),
    .X(_09177_));
 sky130_fd_sc_hd__a22o_1 _15724_ (.A1(\count_instr[41] ),
    .A2(_08802_),
    .B1(_08652_),
    .B2(\count_cycle[41] ),
    .X(_09178_));
 sky130_fd_sc_hd__a221o_1 _15725_ (.A1(\count_instr[9] ),
    .A2(_08749_),
    .B1(\count_cycle[9] ),
    .B2(_08748_),
    .C1(_09178_),
    .X(_09179_));
 sky130_fd_sc_hd__mux2_1 _15726_ (.A0(\cpuregs[18][9] ),
    .A1(\cpuregs[19][9] ),
    .S(_08561_),
    .X(_09180_));
 sky130_fd_sc_hd__buf_2 _15727_ (.A(_08573_),
    .X(_09181_));
 sky130_fd_sc_hd__or2_1 _15728_ (.A(\cpuregs[16][9] ),
    .B(_09181_),
    .X(_09182_));
 sky130_fd_sc_hd__o211a_1 _15729_ (.A1(\cpuregs[17][9] ),
    .A2(_09112_),
    .B1(_08570_),
    .C1(_09182_),
    .X(_09183_));
 sky130_fd_sc_hd__a21oi_1 _15730_ (.A1(_08553_),
    .A2(_09180_),
    .B1(_09183_),
    .Y(_09184_));
 sky130_fd_sc_hd__mux2_1 _15731_ (.A0(\cpuregs[10][9] ),
    .A1(\cpuregs[11][9] ),
    .S(_09083_),
    .X(_09185_));
 sky130_fd_sc_hd__buf_4 _15732_ (.A(_08970_),
    .X(_09186_));
 sky130_fd_sc_hd__mux2_1 _15733_ (.A0(\cpuregs[8][9] ),
    .A1(\cpuregs[9][9] ),
    .S(_09186_),
    .X(_09187_));
 sky130_fd_sc_hd__mux2_1 _15734_ (.A0(_09185_),
    .A1(_09187_),
    .S(_08586_),
    .X(_09188_));
 sky130_fd_sc_hd__mux2_1 _15735_ (.A0(\cpuregs[12][9] ),
    .A1(\cpuregs[13][9] ),
    .S(_08618_),
    .X(_09189_));
 sky130_fd_sc_hd__mux2_1 _15736_ (.A0(\cpuregs[14][9] ),
    .A1(\cpuregs[15][9] ),
    .S(_08595_),
    .X(_09190_));
 sky130_fd_sc_hd__or2_1 _15737_ (.A(_08593_),
    .B(_09190_),
    .X(_09191_));
 sky130_fd_sc_hd__o211a_1 _15738_ (.A1(_09123_),
    .A2(_09189_),
    .B1(_09191_),
    .C1(_08600_),
    .X(_09192_));
 sky130_fd_sc_hd__a211o_1 _15739_ (.A1(_08581_),
    .A2(_09188_),
    .B1(_09192_),
    .C1(_08605_),
    .X(_09193_));
 sky130_fd_sc_hd__mux2_1 _15740_ (.A0(\cpuregs[2][9] ),
    .A1(\cpuregs[3][9] ),
    .S(_09134_),
    .X(_09194_));
 sky130_fd_sc_hd__mux2_1 _15741_ (.A0(\cpuregs[0][9] ),
    .A1(\cpuregs[1][9] ),
    .S(_09136_),
    .X(_09195_));
 sky130_fd_sc_hd__mux2_1 _15742_ (.A0(_09194_),
    .A1(_09195_),
    .S(_08613_),
    .X(_09196_));
 sky130_fd_sc_hd__clkbuf_4 _15743_ (.A(_08970_),
    .X(_09197_));
 sky130_fd_sc_hd__mux2_1 _15744_ (.A0(\cpuregs[4][9] ),
    .A1(\cpuregs[5][9] ),
    .S(_09197_),
    .X(_09198_));
 sky130_fd_sc_hd__mux2_1 _15745_ (.A0(\cpuregs[6][9] ),
    .A1(\cpuregs[7][9] ),
    .S(_08842_),
    .X(_09199_));
 sky130_fd_sc_hd__or2_1 _15746_ (.A(_08735_),
    .B(_09199_),
    .X(_09200_));
 sky130_fd_sc_hd__o211a_1 _15747_ (.A1(_09139_),
    .A2(_09198_),
    .B1(_09200_),
    .C1(_08620_),
    .X(_09201_));
 sky130_fd_sc_hd__buf_2 _15748_ (.A(_08616_),
    .X(_09202_));
 sky130_fd_sc_hd__a211o_1 _15749_ (.A1(_08608_),
    .A2(_09196_),
    .B1(_09201_),
    .C1(_09202_),
    .X(_09203_));
 sky130_fd_sc_hd__a21oi_2 _15750_ (.A1(_09193_),
    .A2(_09203_),
    .B1(_09148_),
    .Y(_09204_));
 sky130_fd_sc_hd__a211o_4 _15751_ (.A1(_08545_),
    .A2(_09184_),
    .B1(_09204_),
    .C1(_09150_),
    .X(_09205_));
 sky130_fd_sc_hd__clkbuf_2 _15752_ (.A(_08936_),
    .X(_09206_));
 sky130_fd_sc_hd__clkbuf_2 _15753_ (.A(_08641_),
    .X(_09207_));
 sky130_fd_sc_hd__a221o_1 _15754_ (.A1(\irq_mask[9] ),
    .A2(_09206_),
    .B1(\timer[9] ),
    .B2(_09207_),
    .C1(_09035_),
    .X(_09208_));
 sky130_fd_sc_hd__o21bai_1 _15755_ (.A1(_08690_),
    .A2(_09205_),
    .B1_N(_09208_),
    .Y(_09209_));
 sky130_fd_sc_hd__buf_2 _15756_ (.A(_08945_),
    .X(_09210_));
 sky130_fd_sc_hd__o211a_1 _15757_ (.A1(_08753_),
    .A2(_09179_),
    .B1(_09209_),
    .C1(_09210_),
    .X(_09211_));
 sky130_fd_sc_hd__mux2_2 _15758_ (.A0(\genblk1.pcpi_mul.rd[9] ),
    .A1(\genblk1.pcpi_mul.rd[41] ),
    .S(_09052_),
    .X(_09212_));
 sky130_fd_sc_hd__buf_2 _15759_ (.A(_08676_),
    .X(_09213_));
 sky130_fd_sc_hd__o221a_1 _15760_ (.A1(net64),
    .A2(_09161_),
    .B1(_09213_),
    .B2(net50),
    .C1(_09164_),
    .X(_09214_));
 sky130_fd_sc_hd__o21a_1 _15761_ (.A1(_09160_),
    .A2(_09214_),
    .B1(_08880_),
    .X(_09215_));
 sky130_fd_sc_hd__a211o_1 _15762_ (.A1(_08902_),
    .A2(_09212_),
    .B1(_09215_),
    .C1(_08666_),
    .X(_09216_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15763_ (.A(_08541_),
    .X(_09217_));
 sky130_fd_sc_hd__o32a_1 _15764_ (.A1(_09177_),
    .A2(_09211_),
    .A3(_09216_),
    .B1(_09217_),
    .B2(\irq_pending[9] ),
    .X(_14603_));
 sky130_fd_sc_hd__clkbuf_2 _15765_ (.A(\reg_pc[10] ),
    .X(_09218_));
 sky130_fd_sc_hd__clkbuf_2 _15766_ (.A(\decoded_imm[10] ),
    .X(_09219_));
 sky130_fd_sc_hd__nor2_1 _15767_ (.A(_09218_),
    .B(_09219_),
    .Y(_09220_));
 sky130_fd_sc_hd__and2_1 _15768_ (.A(\reg_pc[10] ),
    .B(_09219_),
    .X(_09221_));
 sky130_fd_sc_hd__o2111ai_1 _15769_ (.A1(_09220_),
    .A2(_09221_),
    .B1(_09171_),
    .C1(_09175_),
    .D1(_09176_),
    .Y(_09222_));
 sky130_fd_sc_hd__a311o_1 _15770_ (.A1(_09171_),
    .A2(_09175_),
    .A3(_09176_),
    .B1(_09220_),
    .C1(_09221_),
    .X(_09223_));
 sky130_fd_sc_hd__mux2_1 _15771_ (.A0(\cpuregs[18][10] ),
    .A1(\cpuregs[19][10] ),
    .S(_08825_),
    .X(_09224_));
 sky130_fd_sc_hd__or2_1 _15772_ (.A(\cpuregs[16][10] ),
    .B(_08697_),
    .X(_09225_));
 sky130_fd_sc_hd__o211a_1 _15773_ (.A1(\cpuregs[17][10] ),
    .A2(_09055_),
    .B1(_08950_),
    .C1(_09225_),
    .X(_09226_));
 sky130_fd_sc_hd__a21oi_1 _15774_ (.A1(_08948_),
    .A2(_09224_),
    .B1(_09226_),
    .Y(_09227_));
 sky130_fd_sc_hd__mux2_1 _15775_ (.A0(\cpuregs[2][10] ),
    .A1(\cpuregs[3][10] ),
    .S(_09060_),
    .X(_09228_));
 sky130_fd_sc_hd__mux2_1 _15776_ (.A0(\cpuregs[0][10] ),
    .A1(\cpuregs[1][10] ),
    .S(_08833_),
    .X(_09229_));
 sky130_fd_sc_hd__mux2_1 _15777_ (.A0(_09228_),
    .A1(_09229_),
    .S(_08613_),
    .X(_09230_));
 sky130_fd_sc_hd__mux2_1 _15778_ (.A0(\cpuregs[4][10] ),
    .A1(\cpuregs[5][10] ),
    .S(_09066_),
    .X(_09231_));
 sky130_fd_sc_hd__mux2_1 _15779_ (.A0(\cpuregs[6][10] ),
    .A1(\cpuregs[7][10] ),
    .S(_09069_),
    .X(_09232_));
 sky130_fd_sc_hd__or2_1 _15780_ (.A(_09068_),
    .B(_09232_),
    .X(_09233_));
 sky130_fd_sc_hd__o211a_1 _15781_ (.A1(_08839_),
    .A2(_09231_),
    .B1(_09233_),
    .C1(_08845_),
    .X(_09234_));
 sky130_fd_sc_hd__a211o_1 _15782_ (.A1(_08831_),
    .A2(_09230_),
    .B1(_09234_),
    .C1(_09132_),
    .X(_09235_));
 sky130_fd_sc_hd__mux2_1 _15783_ (.A0(\cpuregs[14][10] ),
    .A1(\cpuregs[15][10] ),
    .S(_09076_),
    .X(_09236_));
 sky130_fd_sc_hd__mux2_1 _15784_ (.A0(\cpuregs[12][10] ),
    .A1(\cpuregs[13][10] ),
    .S(_09078_),
    .X(_09237_));
 sky130_fd_sc_hd__mux2_1 _15785_ (.A0(_09236_),
    .A1(_09237_),
    .S(_09018_),
    .X(_09238_));
 sky130_fd_sc_hd__mux2_1 _15786_ (.A0(\cpuregs[8][10] ),
    .A1(\cpuregs[9][10] ),
    .S(_09083_),
    .X(_09239_));
 sky130_fd_sc_hd__mux2_1 _15787_ (.A0(\cpuregs[10][10] ),
    .A1(\cpuregs[11][10] ),
    .S(_08911_),
    .X(_09240_));
 sky130_fd_sc_hd__or2_1 _15788_ (.A(_08730_),
    .B(_09240_),
    .X(_09241_));
 sky130_fd_sc_hd__o211a_1 _15789_ (.A1(_09082_),
    .A2(_09239_),
    .B1(_09241_),
    .C1(_08607_),
    .X(_09242_));
 sky130_fd_sc_hd__a211o_1 _15790_ (.A1(_08860_),
    .A2(_09238_),
    .B1(_09242_),
    .C1(_08975_),
    .X(_09243_));
 sky130_fd_sc_hd__a21oi_2 _15791_ (.A1(_09235_),
    .A2(_09243_),
    .B1(_09090_),
    .Y(_09244_));
 sky130_fd_sc_hd__a211o_4 _15792_ (.A1(_08824_),
    .A2(_09227_),
    .B1(_09244_),
    .C1(_09092_),
    .X(_09245_));
 sky130_fd_sc_hd__nor2_1 _15793_ (.A(_09009_),
    .B(_09245_),
    .Y(_09246_));
 sky130_fd_sc_hd__clkbuf_2 _15794_ (.A(\timer[10] ),
    .X(_09247_));
 sky130_fd_sc_hd__a221o_1 _15795_ (.A1(\irq_mask[10] ),
    .A2(_08638_),
    .B1(_09247_),
    .B2(_08642_),
    .C1(_09035_),
    .X(_09248_));
 sky130_fd_sc_hd__a22o_1 _15796_ (.A1(\count_instr[10] ),
    .A2(_08941_),
    .B1(_08651_),
    .B2(\count_cycle[42] ),
    .X(_09249_));
 sky130_fd_sc_hd__a21o_1 _15797_ (.A1(\count_instr[42] ),
    .A2(_08658_),
    .B1(_09249_),
    .X(_09250_));
 sky130_fd_sc_hd__a211o_1 _15798_ (.A1(\count_cycle[10] ),
    .A2(_09037_),
    .B1(_09250_),
    .C1(_08752_),
    .X(_09251_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15799_ (.A(_08179_),
    .X(_09252_));
 sky130_fd_sc_hd__o211a_1 _15800_ (.A1(_09246_),
    .A2(_09248_),
    .B1(_09251_),
    .C1(_09252_),
    .X(_09253_));
 sky130_fd_sc_hd__mux2_4 _15801_ (.A0(\genblk1.pcpi_mul.rd[10] ),
    .A1(\genblk1.pcpi_mul.rd[42] ),
    .S(_08884_),
    .X(_09254_));
 sky130_fd_sc_hd__o221a_1 _15802_ (.A1(net34),
    .A2(_09161_),
    .B1(_08676_),
    .B2(net51),
    .C1(_09164_),
    .X(_09255_));
 sky130_fd_sc_hd__o21a_1 _15803_ (.A1(_09160_),
    .A2(_09255_),
    .B1(_08152_),
    .X(_09256_));
 sky130_fd_sc_hd__a211o_1 _15804_ (.A1(_08517_),
    .A2(_09254_),
    .B1(_09256_),
    .C1(_08773_),
    .X(_09257_));
 sky130_fd_sc_hd__o22a_1 _15805_ (.A1(\irq_pending[10] ),
    .A2(_09107_),
    .B1(_09253_),
    .B2(_09257_),
    .X(_09258_));
 sky130_fd_sc_hd__a31o_1 _15806_ (.A1(_09101_),
    .A2(_09222_),
    .A3(_09223_),
    .B1(_09258_),
    .X(_14573_));
 sky130_fd_sc_hd__clkbuf_2 _15807_ (.A(_08688_),
    .X(_09259_));
 sky130_fd_sc_hd__mux2_1 _15808_ (.A0(\cpuregs[16][11] ),
    .A1(\cpuregs[17][11] ),
    .S(_08561_),
    .X(_09260_));
 sky130_fd_sc_hd__or2_1 _15809_ (.A(\cpuregs[18][11] ),
    .B(_08574_),
    .X(_09261_));
 sky130_fd_sc_hd__o211a_1 _15810_ (.A1(\cpuregs[19][11] ),
    .A2(_08565_),
    .B1(_08552_),
    .C1(_09261_),
    .X(_09262_));
 sky130_fd_sc_hd__a21oi_1 _15811_ (.A1(_08702_),
    .A2(_09260_),
    .B1(_09262_),
    .Y(_09263_));
 sky130_fd_sc_hd__buf_4 _15812_ (.A(_08694_),
    .X(_09264_));
 sky130_fd_sc_hd__mux2_1 _15813_ (.A0(\cpuregs[6][11] ),
    .A1(\cpuregs[7][11] ),
    .S(_09264_),
    .X(_09265_));
 sky130_fd_sc_hd__mux2_1 _15814_ (.A0(\cpuregs[4][11] ),
    .A1(\cpuregs[5][11] ),
    .S(_09264_),
    .X(_09266_));
 sky130_fd_sc_hd__mux2_1 _15815_ (.A0(_09265_),
    .A1(_09266_),
    .S(_09018_),
    .X(_09267_));
 sky130_fd_sc_hd__mux2_1 _15816_ (.A0(\cpuregs[2][11] ),
    .A1(\cpuregs[3][11] ),
    .S(_08840_),
    .X(_09268_));
 sky130_fd_sc_hd__or2_1 _15817_ (.A(_08736_),
    .B(_09268_),
    .X(_09269_));
 sky130_fd_sc_hd__mux2_1 _15818_ (.A0(\cpuregs[0][11] ),
    .A1(\cpuregs[1][11] ),
    .S(_08590_),
    .X(_09270_));
 sky130_fd_sc_hd__o21a_1 _15819_ (.A1(_08551_),
    .A2(_09270_),
    .B1(_08580_),
    .X(_09271_));
 sky130_fd_sc_hd__a221o_1 _15820_ (.A1(_08860_),
    .A2(_09267_),
    .B1(_09269_),
    .B2(_09271_),
    .C1(_09202_),
    .X(_09272_));
 sky130_fd_sc_hd__mux2_1 _15821_ (.A0(\cpuregs[8][11] ),
    .A1(\cpuregs[9][11] ),
    .S(_09062_),
    .X(_09273_));
 sky130_fd_sc_hd__mux2_1 _15822_ (.A0(\cpuregs[10][11] ),
    .A1(\cpuregs[11][11] ),
    .S(_08833_),
    .X(_09274_));
 sky130_fd_sc_hd__mux2_1 _15823_ (.A0(_09273_),
    .A1(_09274_),
    .S(_08837_),
    .X(_09275_));
 sky130_fd_sc_hd__mux2_1 _15824_ (.A0(\cpuregs[12][11] ),
    .A1(\cpuregs[13][11] ),
    .S(_09066_),
    .X(_09276_));
 sky130_fd_sc_hd__mux2_1 _15825_ (.A0(\cpuregs[14][11] ),
    .A1(\cpuregs[15][11] ),
    .S(_08842_),
    .X(_09277_));
 sky130_fd_sc_hd__or2_1 _15826_ (.A(_08735_),
    .B(_09277_),
    .X(_09278_));
 sky130_fd_sc_hd__o211a_1 _15827_ (.A1(_08839_),
    .A2(_09276_),
    .B1(_09278_),
    .C1(_08845_),
    .X(_09279_));
 sky130_fd_sc_hd__a211o_1 _15828_ (.A1(_08831_),
    .A2(_09275_),
    .B1(_09279_),
    .C1(_09073_),
    .X(_09280_));
 sky130_fd_sc_hd__a21oi_2 _15829_ (.A1(_09272_),
    .A2(_09280_),
    .B1(_08627_),
    .Y(_09281_));
 sky130_fd_sc_hd__a211o_4 _15830_ (.A1(_08545_),
    .A2(_09263_),
    .B1(_09281_),
    .C1(_08634_),
    .X(_09282_));
 sky130_fd_sc_hd__nor2_1 _15831_ (.A(_09259_),
    .B(_09282_),
    .Y(_09283_));
 sky130_fd_sc_hd__a221o_1 _15832_ (.A1(\irq_mask[11] ),
    .A2(_09206_),
    .B1(\timer[11] ),
    .B2(_08642_),
    .C1(_09035_),
    .X(_09284_));
 sky130_fd_sc_hd__clkbuf_2 _15833_ (.A(_08656_),
    .X(_09285_));
 sky130_fd_sc_hd__clkbuf_2 _15834_ (.A(_08804_),
    .X(_09286_));
 sky130_fd_sc_hd__a22o_1 _15835_ (.A1(\count_instr[43] ),
    .A2(_08942_),
    .B1(_09286_),
    .B2(\count_cycle[43] ),
    .X(_09287_));
 sky130_fd_sc_hd__a221o_1 _15836_ (.A1(\count_instr[11] ),
    .A2(_09285_),
    .B1(\count_cycle[11] ),
    .B2(_08654_),
    .C1(_09287_),
    .X(_09288_));
 sky130_fd_sc_hd__o22a_1 _15837_ (.A1(_09283_),
    .A2(_09284_),
    .B1(_09288_),
    .B2(_08650_),
    .X(_09289_));
 sky130_fd_sc_hd__mux2_2 _15838_ (.A0(\genblk1.pcpi_mul.rd[11] ),
    .A1(\genblk1.pcpi_mul.rd[43] ),
    .S(_08900_),
    .X(_09290_));
 sky130_fd_sc_hd__clkbuf_2 _15839_ (.A(_08517_),
    .X(_09291_));
 sky130_fd_sc_hd__a22o_1 _15840_ (.A1(_09210_),
    .A2(_09289_),
    .B1(_09290_),
    .B2(_09291_),
    .X(_09292_));
 sky130_fd_sc_hd__nand2_1 _15841_ (.A(_09218_),
    .B(_09219_),
    .Y(_09293_));
 sky130_fd_sc_hd__or2_1 _15842_ (.A(\reg_pc[11] ),
    .B(\decoded_imm[11] ),
    .X(_09294_));
 sky130_fd_sc_hd__clkbuf_2 _15843_ (.A(\reg_pc[11] ),
    .X(_09295_));
 sky130_fd_sc_hd__nand2_1 _15844_ (.A(_09295_),
    .B(\decoded_imm[11] ),
    .Y(_09296_));
 sky130_fd_sc_hd__nand2_1 _15845_ (.A(_09294_),
    .B(_09296_),
    .Y(_09297_));
 sky130_fd_sc_hd__a21oi_2 _15846_ (.A1(_09293_),
    .A2(_09223_),
    .B1(_09297_),
    .Y(_09298_));
 sky130_fd_sc_hd__clkbuf_4 _15847_ (.A(_08295_),
    .X(_09299_));
 sky130_fd_sc_hd__a31o_1 _15848_ (.A1(_09293_),
    .A2(_09223_),
    .A3(_09297_),
    .B1(_09299_),
    .X(_09300_));
 sky130_fd_sc_hd__o221a_1 _15849_ (.A1(net35),
    .A2(_09161_),
    .B1(_09213_),
    .B2(net52),
    .C1(_09164_),
    .X(_09301_));
 sky130_fd_sc_hd__o21ai_1 _15850_ (.A1(_09160_),
    .A2(_09301_),
    .B1(_08231_),
    .Y(_09302_));
 sky130_fd_sc_hd__o211ai_1 _15851_ (.A1(_09298_),
    .A2(_09300_),
    .B1(_09302_),
    .C1(_08541_),
    .Y(_09303_));
 sky130_fd_sc_hd__o22a_1 _15852_ (.A1(\irq_pending[11] ),
    .A2(_09217_),
    .B1(_09292_),
    .B2(_09303_),
    .X(_14574_));
 sky130_vsdinv _15853_ (.A(_09296_),
    .Y(_09304_));
 sky130_fd_sc_hd__clkbuf_2 _15854_ (.A(\decoded_imm[12] ),
    .X(_09305_));
 sky130_fd_sc_hd__or2_1 _15855_ (.A(\reg_pc[12] ),
    .B(_09305_),
    .X(_09306_));
 sky130_fd_sc_hd__nand2_2 _15856_ (.A(\reg_pc[12] ),
    .B(_09305_),
    .Y(_09307_));
 sky130_fd_sc_hd__o211a_1 _15857_ (.A1(_09304_),
    .A2(_09298_),
    .B1(_09306_),
    .C1(_09307_),
    .X(_09308_));
 sky130_fd_sc_hd__a211o_1 _15858_ (.A1(_09306_),
    .A2(_09307_),
    .B1(_09304_),
    .C1(_09298_),
    .X(_09309_));
 sky130_fd_sc_hd__and3b_1 _15859_ (.A_N(_09308_),
    .B(_09309_),
    .C(_08894_),
    .X(_09310_));
 sky130_fd_sc_hd__mux2_1 _15860_ (.A0(\cpuregs[16][12] ),
    .A1(\cpuregs[17][12] ),
    .S(_08825_),
    .X(_09311_));
 sky130_fd_sc_hd__or2_1 _15861_ (.A(\cpuregs[18][12] ),
    .B(_08697_),
    .X(_09312_));
 sky130_fd_sc_hd__o211a_1 _15862_ (.A1(\cpuregs[19][12] ),
    .A2(_09055_),
    .B1(_08716_),
    .C1(_09312_),
    .X(_09313_));
 sky130_fd_sc_hd__a21oi_1 _15863_ (.A1(_08701_),
    .A2(_09311_),
    .B1(_09313_),
    .Y(_09314_));
 sky130_fd_sc_hd__mux2_1 _15864_ (.A0(\cpuregs[6][12] ),
    .A1(\cpuregs[7][12] ),
    .S(_08610_),
    .X(_09315_));
 sky130_fd_sc_hd__or2_1 _15865_ (.A(_08731_),
    .B(_09315_),
    .X(_09316_));
 sky130_fd_sc_hd__mux2_1 _15866_ (.A0(\cpuregs[4][12] ),
    .A1(\cpuregs[5][12] ),
    .S(_08582_),
    .X(_09317_));
 sky130_fd_sc_hd__o21a_1 _15867_ (.A1(_08839_),
    .A2(_09317_),
    .B1(_08859_),
    .X(_09318_));
 sky130_fd_sc_hd__mux2_1 _15868_ (.A0(\cpuregs[2][12] ),
    .A1(\cpuregs[3][12] ),
    .S(_09078_),
    .X(_09319_));
 sky130_fd_sc_hd__mux2_1 _15869_ (.A0(\cpuregs[0][12] ),
    .A1(\cpuregs[1][12] ),
    .S(_09264_),
    .X(_09320_));
 sky130_fd_sc_hd__mux2_1 _15870_ (.A0(_09319_),
    .A1(_09320_),
    .S(_09018_),
    .X(_09321_));
 sky130_fd_sc_hd__a221o_1 _15871_ (.A1(_09316_),
    .A2(_09318_),
    .B1(_09321_),
    .B2(_08954_),
    .C1(_08617_),
    .X(_09322_));
 sky130_fd_sc_hd__mux2_1 _15872_ (.A0(\cpuregs[8][12] ),
    .A1(\cpuregs[9][12] ),
    .S(_09076_),
    .X(_09323_));
 sky130_fd_sc_hd__mux2_1 _15873_ (.A0(\cpuregs[10][12] ),
    .A1(\cpuregs[11][12] ),
    .S(_09078_),
    .X(_09324_));
 sky130_fd_sc_hd__mux2_1 _15874_ (.A0(_09323_),
    .A1(_09324_),
    .S(_08967_),
    .X(_09325_));
 sky130_fd_sc_hd__mux2_1 _15875_ (.A0(\cpuregs[12][12] ),
    .A1(\cpuregs[13][12] ),
    .S(_09083_),
    .X(_09326_));
 sky130_fd_sc_hd__mux2_1 _15876_ (.A0(\cpuregs[14][12] ),
    .A1(\cpuregs[15][12] ),
    .S(_08911_),
    .X(_09327_));
 sky130_fd_sc_hd__or2_1 _15877_ (.A(_08730_),
    .B(_09327_),
    .X(_09328_));
 sky130_fd_sc_hd__o211a_1 _15878_ (.A1(_09082_),
    .A2(_09326_),
    .B1(_09328_),
    .C1(_09087_),
    .X(_09329_));
 sky130_fd_sc_hd__a211o_1 _15879_ (.A1(_09075_),
    .A2(_09325_),
    .B1(_09329_),
    .C1(_08975_),
    .X(_09330_));
 sky130_fd_sc_hd__a21oi_2 _15880_ (.A1(_09322_),
    .A2(_09330_),
    .B1(_09090_),
    .Y(_09331_));
 sky130_fd_sc_hd__a211o_4 _15881_ (.A1(_08824_),
    .A2(_09314_),
    .B1(_09331_),
    .C1(_09092_),
    .X(_09332_));
 sky130_fd_sc_hd__nor2_1 _15882_ (.A(_08689_),
    .B(_09332_),
    .Y(_09333_));
 sky130_fd_sc_hd__a221o_1 _15883_ (.A1(\irq_mask[12] ),
    .A2(_08937_),
    .B1(\timer[12] ),
    .B2(_08938_),
    .C1(_08939_),
    .X(_09334_));
 sky130_fd_sc_hd__a22o_1 _15884_ (.A1(\count_instr[44] ),
    .A2(_08801_),
    .B1(_08651_),
    .B2(\count_cycle[44] ),
    .X(_09335_));
 sky130_fd_sc_hd__a221o_1 _15885_ (.A1(\count_instr[12] ),
    .A2(_08803_),
    .B1(\count_cycle[12] ),
    .B2(_08747_),
    .C1(_09335_),
    .X(_09336_));
 sky130_fd_sc_hd__clkbuf_2 _15886_ (.A(_08649_),
    .X(_09337_));
 sky130_fd_sc_hd__o22a_1 _15887_ (.A1(_09333_),
    .A2(_09334_),
    .B1(_09336_),
    .B2(_09337_),
    .X(_09338_));
 sky130_fd_sc_hd__mux2_4 _15888_ (.A0(\genblk1.pcpi_mul.rd[12] ),
    .A1(\genblk1.pcpi_mul.rd[44] ),
    .S(_09052_),
    .X(_09339_));
 sky130_fd_sc_hd__o221a_1 _15889_ (.A1(net36),
    .A2(_09161_),
    .B1(_09213_),
    .B2(net53),
    .C1(_09164_),
    .X(_09340_));
 sky130_fd_sc_hd__o21a_1 _15890_ (.A1(_09160_),
    .A2(_09340_),
    .B1(_08230_),
    .X(_09341_));
 sky130_fd_sc_hd__a221o_1 _15891_ (.A1(_08180_),
    .A2(_09338_),
    .B1(_09339_),
    .B2(_08902_),
    .C1(_09341_),
    .X(_09342_));
 sky130_fd_sc_hd__a211o_1 _15892_ (.A1(\irq_pending[12] ),
    .A2(_08774_),
    .B1(_09310_),
    .C1(_09342_),
    .X(_14575_));
 sky130_fd_sc_hd__and2_1 _15893_ (.A(\reg_pc[13] ),
    .B(\decoded_imm[13] ),
    .X(_09343_));
 sky130_fd_sc_hd__nor2_1 _15894_ (.A(\reg_pc[13] ),
    .B(\decoded_imm[13] ),
    .Y(_09344_));
 sky130_fd_sc_hd__nor2_1 _15895_ (.A(_09343_),
    .B(_09344_),
    .Y(_09345_));
 sky130_fd_sc_hd__o2111ai_2 _15896_ (.A1(_09304_),
    .A2(_09298_),
    .B1(_09306_),
    .C1(_09307_),
    .D1(_09345_),
    .Y(_09346_));
 sky130_fd_sc_hd__clkbuf_2 _15897_ (.A(\reg_pc[12] ),
    .X(_09347_));
 sky130_fd_sc_hd__a21o_1 _15898_ (.A1(_09347_),
    .A2(_09305_),
    .B1(_09308_),
    .X(_09348_));
 sky130_fd_sc_hd__mux2_1 _15899_ (.A0(_09348_),
    .A1(_09307_),
    .S(_09345_),
    .X(_09349_));
 sky130_fd_sc_hd__and3_1 _15900_ (.A(_08894_),
    .B(_09346_),
    .C(_09349_),
    .X(_09350_));
 sky130_fd_sc_hd__mux2_1 _15901_ (.A0(\cpuregs[16][13] ),
    .A1(\cpuregs[17][13] ),
    .S(_08825_),
    .X(_09351_));
 sky130_fd_sc_hd__or2_1 _15902_ (.A(\cpuregs[18][13] ),
    .B(_08697_),
    .X(_09352_));
 sky130_fd_sc_hd__o211a_1 _15903_ (.A1(\cpuregs[19][13] ),
    .A2(_08827_),
    .B1(_08716_),
    .C1(_09352_),
    .X(_09353_));
 sky130_fd_sc_hd__a21oi_1 _15904_ (.A1(_08701_),
    .A2(_09351_),
    .B1(_09353_),
    .Y(_09354_));
 sky130_fd_sc_hd__mux2_1 _15905_ (.A0(\cpuregs[8][13] ),
    .A1(\cpuregs[9][13] ),
    .S(_09060_),
    .X(_09355_));
 sky130_fd_sc_hd__mux2_1 _15906_ (.A0(\cpuregs[10][13] ),
    .A1(\cpuregs[11][13] ),
    .S(_08833_),
    .X(_09356_));
 sky130_fd_sc_hd__mux2_1 _15907_ (.A0(_09355_),
    .A1(_09356_),
    .S(_08837_),
    .X(_09357_));
 sky130_fd_sc_hd__mux2_1 _15908_ (.A0(\cpuregs[12][13] ),
    .A1(\cpuregs[13][13] ),
    .S(_09066_),
    .X(_09358_));
 sky130_fd_sc_hd__mux2_1 _15909_ (.A0(\cpuregs[14][13] ),
    .A1(\cpuregs[15][13] ),
    .S(_09069_),
    .X(_09359_));
 sky130_fd_sc_hd__or2_1 _15910_ (.A(_09068_),
    .B(_09359_),
    .X(_09360_));
 sky130_fd_sc_hd__o211a_1 _15911_ (.A1(_08839_),
    .A2(_09358_),
    .B1(_09360_),
    .C1(_08845_),
    .X(_09361_));
 sky130_fd_sc_hd__a211o_1 _15912_ (.A1(_08831_),
    .A2(_09357_),
    .B1(_09361_),
    .C1(_09073_),
    .X(_09362_));
 sky130_fd_sc_hd__mux2_1 _15913_ (.A0(\cpuregs[2][13] ),
    .A1(\cpuregs[3][13] ),
    .S(_09264_),
    .X(_09363_));
 sky130_fd_sc_hd__or2_1 _15914_ (.A(_08731_),
    .B(_09363_),
    .X(_09364_));
 sky130_fd_sc_hd__mux2_1 _15915_ (.A0(\cpuregs[0][13] ),
    .A1(\cpuregs[1][13] ),
    .S(_08835_),
    .X(_09365_));
 sky130_fd_sc_hd__o21a_1 _15916_ (.A1(_08851_),
    .A2(_09365_),
    .B1(_08706_),
    .X(_09366_));
 sky130_fd_sc_hd__mux2_1 _15917_ (.A0(\cpuregs[6][13] ),
    .A1(\cpuregs[7][13] ),
    .S(_08559_),
    .X(_09367_));
 sky130_fd_sc_hd__mux2_1 _15918_ (.A0(\cpuregs[4][13] ),
    .A1(\cpuregs[5][13] ),
    .S(_08559_),
    .X(_09368_));
 sky130_fd_sc_hd__mux2_1 _15919_ (.A0(_09367_),
    .A1(_09368_),
    .S(_08857_),
    .X(_09369_));
 sky130_fd_sc_hd__a221o_1 _15920_ (.A1(_09364_),
    .A2(_09366_),
    .B1(_09369_),
    .B2(_08860_),
    .C1(_08861_),
    .X(_09370_));
 sky130_fd_sc_hd__a21oi_1 _15921_ (.A1(_09362_),
    .A2(_09370_),
    .B1(_08691_),
    .Y(_09371_));
 sky130_fd_sc_hd__a211o_4 _15922_ (.A1(_08824_),
    .A2(_09354_),
    .B1(_09371_),
    .C1(_08864_),
    .X(_09372_));
 sky130_fd_sc_hd__nor2_1 _15923_ (.A(_09259_),
    .B(_09372_),
    .Y(_09373_));
 sky130_fd_sc_hd__a221o_1 _15924_ (.A1(\irq_mask[13] ),
    .A2(_08638_),
    .B1(\timer[13] ),
    .B2(_08642_),
    .C1(_09035_),
    .X(_09374_));
 sky130_fd_sc_hd__clkbuf_2 _15925_ (.A(_08657_),
    .X(_09375_));
 sky130_fd_sc_hd__a22o_1 _15926_ (.A1(\count_instr[45] ),
    .A2(_09375_),
    .B1(_09286_),
    .B2(\count_cycle[45] ),
    .X(_09376_));
 sky130_fd_sc_hd__a221o_1 _15927_ (.A1(\count_instr[13] ),
    .A2(_09285_),
    .B1(\count_cycle[13] ),
    .B2(_08654_),
    .C1(_09376_),
    .X(_09377_));
 sky130_fd_sc_hd__clkbuf_2 _15928_ (.A(_08649_),
    .X(_09378_));
 sky130_fd_sc_hd__o22a_1 _15929_ (.A1(_09373_),
    .A2(_09374_),
    .B1(_09377_),
    .B2(_09378_),
    .X(_09379_));
 sky130_fd_sc_hd__o221a_1 _15930_ (.A1(net37),
    .A2(_08674_),
    .B1(_08676_),
    .B2(net54),
    .C1(_09163_),
    .X(_09380_));
 sky130_fd_sc_hd__or2_1 _15931_ (.A(_09159_),
    .B(_09380_),
    .X(_09381_));
 sky130_fd_sc_hd__mux2_2 _15932_ (.A0(\genblk1.pcpi_mul.rd[13] ),
    .A1(\genblk1.pcpi_mul.rd[45] ),
    .S(_08884_),
    .X(_09382_));
 sky130_fd_sc_hd__a22o_1 _15933_ (.A1(_08880_),
    .A2(_09381_),
    .B1(_09382_),
    .B2(_08886_),
    .X(_09383_));
 sky130_fd_sc_hd__a211o_1 _15934_ (.A1(_09210_),
    .A2(_09379_),
    .B1(_09383_),
    .C1(_08810_),
    .X(_09384_));
 sky130_fd_sc_hd__o22a_1 _15935_ (.A1(\irq_pending[13] ),
    .A2(_09217_),
    .B1(_09350_),
    .B2(_09384_),
    .X(_14576_));
 sky130_fd_sc_hd__or2_1 _15936_ (.A(\reg_pc[14] ),
    .B(\decoded_imm[14] ),
    .X(_09385_));
 sky130_fd_sc_hd__clkbuf_2 _15937_ (.A(\reg_pc[14] ),
    .X(_09386_));
 sky130_fd_sc_hd__nand2_1 _15938_ (.A(_09386_),
    .B(\decoded_imm[14] ),
    .Y(_09387_));
 sky130_fd_sc_hd__nand2_1 _15939_ (.A(_09385_),
    .B(_09387_),
    .Y(_09388_));
 sky130_fd_sc_hd__o21ba_1 _15940_ (.A1(_09307_),
    .A2(_09344_),
    .B1_N(_09343_),
    .X(_09389_));
 sky130_fd_sc_hd__a31o_1 _15941_ (.A1(_09346_),
    .A2(_09388_),
    .A3(_09389_),
    .B1(_08295_),
    .X(_09390_));
 sky130_fd_sc_hd__a21o_1 _15942_ (.A1(_09346_),
    .A2(_09389_),
    .B1(_09388_),
    .X(_09391_));
 sky130_fd_sc_hd__and2b_1 _15943_ (.A_N(_09390_),
    .B(_09391_),
    .X(_09392_));
 sky130_fd_sc_hd__mux2_1 _15944_ (.A0(\cpuregs[18][14] ),
    .A1(\cpuregs[19][14] ),
    .S(_08698_),
    .X(_09393_));
 sky130_fd_sc_hd__or2_1 _15945_ (.A(\cpuregs[16][14] ),
    .B(_08825_),
    .X(_09394_));
 sky130_fd_sc_hd__o211a_1 _15946_ (.A1(\cpuregs[17][14] ),
    .A2(_08700_),
    .B1(_08701_),
    .C1(_09394_),
    .X(_09395_));
 sky130_fd_sc_hd__a21oi_1 _15947_ (.A1(_08693_),
    .A2(_09393_),
    .B1(_09395_),
    .Y(_09396_));
 sky130_fd_sc_hd__mux2_1 _15948_ (.A0(\cpuregs[10][14] ),
    .A1(\cpuregs[11][14] ),
    .S(_08909_),
    .X(_09397_));
 sky130_fd_sc_hd__mux2_1 _15949_ (.A0(\cpuregs[8][14] ),
    .A1(\cpuregs[9][14] ),
    .S(_08909_),
    .X(_09398_));
 sky130_fd_sc_hd__mux2_1 _15950_ (.A0(_09397_),
    .A1(_09398_),
    .S(_08569_),
    .X(_09399_));
 sky130_fd_sc_hd__mux2_1 _15951_ (.A0(\cpuregs[12][14] ),
    .A1(\cpuregs[13][14] ),
    .S(_08696_),
    .X(_09400_));
 sky130_fd_sc_hd__mux2_1 _15952_ (.A0(\cpuregs[14][14] ),
    .A1(\cpuregs[15][14] ),
    .S(_08918_),
    .X(_09401_));
 sky130_fd_sc_hd__or2_1 _15953_ (.A(_08917_),
    .B(_09401_),
    .X(_09402_));
 sky130_fd_sc_hd__o211a_1 _15954_ (.A1(_08915_),
    .A2(_09400_),
    .B1(_09402_),
    .C1(_08921_),
    .X(_09403_));
 sky130_fd_sc_hd__a211o_1 _15955_ (.A1(_08708_),
    .A2(_09399_),
    .B1(_09403_),
    .C1(_08726_),
    .X(_09404_));
 sky130_fd_sc_hd__mux2_1 _15956_ (.A0(\cpuregs[2][14] ),
    .A1(\cpuregs[3][14] ),
    .S(_08912_),
    .X(_09405_));
 sky130_fd_sc_hd__mux2_1 _15957_ (.A0(\cpuregs[0][14] ),
    .A1(\cpuregs[1][14] ),
    .S(_08912_),
    .X(_09406_));
 sky130_fd_sc_hd__mux2_1 _15958_ (.A0(_09405_),
    .A1(_09406_),
    .S(_08721_),
    .X(_09407_));
 sky130_fd_sc_hd__mux2_1 _15959_ (.A0(\cpuregs[4][14] ),
    .A1(\cpuregs[5][14] ),
    .S(_08909_),
    .X(_09408_));
 sky130_fd_sc_hd__mux2_1 _15960_ (.A0(\cpuregs[6][14] ),
    .A1(\cpuregs[7][14] ),
    .S(_08717_),
    .X(_09409_));
 sky130_fd_sc_hd__or2_1 _15961_ (.A(_08917_),
    .B(_09409_),
    .X(_09410_));
 sky130_fd_sc_hd__o211a_1 _15962_ (.A1(_08915_),
    .A2(_09408_),
    .B1(_09410_),
    .C1(_08921_),
    .X(_09411_));
 sky130_fd_sc_hd__a211o_1 _15963_ (.A1(_08708_),
    .A2(_09407_),
    .B1(_09411_),
    .C1(_08740_),
    .X(_09412_));
 sky130_fd_sc_hd__a21oi_1 _15964_ (.A1(_09404_),
    .A2(_09412_),
    .B1(_08824_),
    .Y(_09413_));
 sky130_fd_sc_hd__a211o_4 _15965_ (.A1(_08692_),
    .A2(_09396_),
    .B1(_09413_),
    .C1(_08743_),
    .X(_09414_));
 sky130_fd_sc_hd__nor2_1 _15966_ (.A(_08689_),
    .B(_09414_),
    .Y(_09415_));
 sky130_fd_sc_hd__a221o_1 _15967_ (.A1(\irq_mask[14] ),
    .A2(_08937_),
    .B1(\timer[14] ),
    .B2(_08938_),
    .C1(_09095_),
    .X(_09416_));
 sky130_fd_sc_hd__a22o_1 _15968_ (.A1(\count_instr[46] ),
    .A2(_08801_),
    .B1(_08651_),
    .B2(\count_cycle[46] ),
    .X(_09417_));
 sky130_fd_sc_hd__a221o_1 _15969_ (.A1(\count_instr[14] ),
    .A2(_08803_),
    .B1(\count_cycle[14] ),
    .B2(_08747_),
    .C1(_09417_),
    .X(_09418_));
 sky130_fd_sc_hd__o22a_1 _15970_ (.A1(_09415_),
    .A2(_09416_),
    .B1(_09418_),
    .B2(_09337_),
    .X(_09419_));
 sky130_fd_sc_hd__mux2_4 _15971_ (.A0(\genblk1.pcpi_mul.rd[14] ),
    .A1(\genblk1.pcpi_mul.rd[46] ),
    .S(_09052_),
    .X(_09420_));
 sky130_fd_sc_hd__o221a_1 _15972_ (.A1(net38),
    .A2(_09161_),
    .B1(_09213_),
    .B2(net56),
    .C1(_09164_),
    .X(_09421_));
 sky130_fd_sc_hd__o21a_1 _15973_ (.A1(_09160_),
    .A2(_09421_),
    .B1(_08230_),
    .X(_09422_));
 sky130_fd_sc_hd__a221o_1 _15974_ (.A1(_08180_),
    .A2(_09419_),
    .B1(_09420_),
    .B2(_08902_),
    .C1(_09422_),
    .X(_09423_));
 sky130_fd_sc_hd__a211o_1 _15975_ (.A1(\irq_pending[14] ),
    .A2(_08774_),
    .B1(_09392_),
    .C1(_09423_),
    .X(_14577_));
 sky130_fd_sc_hd__and2_1 _15976_ (.A(\reg_pc[15] ),
    .B(\decoded_imm[15] ),
    .X(_09424_));
 sky130_fd_sc_hd__nor2_1 _15977_ (.A(\reg_pc[15] ),
    .B(\decoded_imm[15] ),
    .Y(_09425_));
 sky130_fd_sc_hd__or2_1 _15978_ (.A(_09424_),
    .B(_09425_),
    .X(_09426_));
 sky130_fd_sc_hd__and2_1 _15979_ (.A(_09387_),
    .B(_09391_),
    .X(_09427_));
 sky130_fd_sc_hd__o21ai_1 _15980_ (.A1(_09426_),
    .A2(_09427_),
    .B1(_08872_),
    .Y(_09428_));
 sky130_fd_sc_hd__a21oi_1 _15981_ (.A1(_09426_),
    .A2(_09427_),
    .B1(_09428_),
    .Y(_09429_));
 sky130_fd_sc_hd__a22o_1 _15982_ (.A1(\count_instr[47] ),
    .A2(_08802_),
    .B1(_08652_),
    .B2(\count_cycle[47] ),
    .X(_09430_));
 sky130_fd_sc_hd__a221o_1 _15983_ (.A1(\count_instr[15] ),
    .A2(_08749_),
    .B1(\count_cycle[15] ),
    .B2(_08748_),
    .C1(_09430_),
    .X(_09431_));
 sky130_fd_sc_hd__mux2_1 _15984_ (.A0(\cpuregs[16][15] ),
    .A1(\cpuregs[17][15] ),
    .S(_08904_),
    .X(_09432_));
 sky130_fd_sc_hd__or2_1 _15985_ (.A(\cpuregs[18][15] ),
    .B(_08574_),
    .X(_09433_));
 sky130_fd_sc_hd__o211a_1 _15986_ (.A1(\cpuregs[19][15] ),
    .A2(_08565_),
    .B1(_08552_),
    .C1(_09433_),
    .X(_09434_));
 sky130_fd_sc_hd__a21oi_1 _15987_ (.A1(_08702_),
    .A2(_09432_),
    .B1(_09434_),
    .Y(_09435_));
 sky130_fd_sc_hd__mux2_1 _15988_ (.A0(\cpuregs[6][15] ),
    .A1(\cpuregs[7][15] ),
    .S(_08582_),
    .X(_09436_));
 sky130_fd_sc_hd__or2_1 _15989_ (.A(_08736_),
    .B(_09436_),
    .X(_09437_));
 sky130_fd_sc_hd__mux2_1 _15990_ (.A0(\cpuregs[4][15] ),
    .A1(\cpuregs[5][15] ),
    .S(_08590_),
    .X(_09438_));
 sky130_fd_sc_hd__o21a_1 _15991_ (.A1(_08589_),
    .A2(_09438_),
    .B1(_08845_),
    .X(_09439_));
 sky130_fd_sc_hd__mux2_1 _15992_ (.A0(\cpuregs[2][15] ),
    .A1(\cpuregs[3][15] ),
    .S(_08833_),
    .X(_09440_));
 sky130_fd_sc_hd__mux2_1 _15993_ (.A0(\cpuregs[0][15] ),
    .A1(\cpuregs[1][15] ),
    .S(_08835_),
    .X(_09441_));
 sky130_fd_sc_hd__mux2_1 _15994_ (.A0(_09440_),
    .A1(_09441_),
    .S(_08613_),
    .X(_09442_));
 sky130_fd_sc_hd__a221o_1 _15995_ (.A1(_09437_),
    .A2(_09439_),
    .B1(_09442_),
    .B2(_09075_),
    .C1(_09202_),
    .X(_09443_));
 sky130_fd_sc_hd__mux2_1 _15996_ (.A0(\cpuregs[8][15] ),
    .A1(\cpuregs[9][15] ),
    .S(_09118_),
    .X(_09444_));
 sky130_fd_sc_hd__mux2_1 _15997_ (.A0(\cpuregs[10][15] ),
    .A1(\cpuregs[11][15] ),
    .S(_09062_),
    .X(_09445_));
 sky130_fd_sc_hd__mux2_1 _15998_ (.A0(_09444_),
    .A1(_09445_),
    .S(_08851_),
    .X(_09446_));
 sky130_fd_sc_hd__mux2_1 _15999_ (.A0(\cpuregs[12][15] ),
    .A1(\cpuregs[13][15] ),
    .S(_09124_),
    .X(_09447_));
 sky130_fd_sc_hd__mux2_1 _16000_ (.A0(\cpuregs[14][15] ),
    .A1(\cpuregs[15][15] ),
    .S(_09127_),
    .X(_09448_));
 sky130_fd_sc_hd__or2_1 _16001_ (.A(_09126_),
    .B(_09448_),
    .X(_09449_));
 sky130_fd_sc_hd__o211a_1 _16002_ (.A1(_09065_),
    .A2(_09447_),
    .B1(_09449_),
    .C1(_09130_),
    .X(_09450_));
 sky130_fd_sc_hd__a211o_1 _16003_ (.A1(_09117_),
    .A2(_09446_),
    .B1(_09450_),
    .C1(_08605_),
    .X(_09451_));
 sky130_fd_sc_hd__a21oi_2 _16004_ (.A1(_09443_),
    .A2(_09451_),
    .B1(_08627_),
    .Y(_09452_));
 sky130_fd_sc_hd__a211o_4 _16005_ (.A1(_08903_),
    .A2(_09435_),
    .B1(_09452_),
    .C1(_08634_),
    .X(_09453_));
 sky130_fd_sc_hd__a221o_1 _16006_ (.A1(\irq_mask[15] ),
    .A2(_09206_),
    .B1(\timer[15] ),
    .B2(_09207_),
    .C1(_09035_),
    .X(_09454_));
 sky130_fd_sc_hd__o21bai_1 _16007_ (.A1(_08690_),
    .A2(_09453_),
    .B1_N(_09454_),
    .Y(_09455_));
 sky130_fd_sc_hd__o211a_1 _16008_ (.A1(_08753_),
    .A2(_09431_),
    .B1(_09455_),
    .C1(_09210_),
    .X(_09456_));
 sky130_fd_sc_hd__mux2_2 _16009_ (.A0(\genblk1.pcpi_mul.rd[15] ),
    .A1(\genblk1.pcpi_mul.rd[47] ),
    .S(_09052_),
    .X(_09457_));
 sky130_fd_sc_hd__a21o_1 _16010_ (.A1(_08324_),
    .A2(_09049_),
    .B1(_08673_),
    .X(_09458_));
 sky130_fd_sc_hd__o21a_1 _16011_ (.A1(net39),
    .A2(_08674_),
    .B1(_09458_),
    .X(_09459_));
 sky130_fd_sc_hd__or2_1 _16012_ (.A(latched_is_lb),
    .B(latched_is_lh),
    .X(_09460_));
 sky130_fd_sc_hd__clkbuf_2 _16013_ (.A(_09460_),
    .X(_09461_));
 sky130_vsdinv _16014_ (.A(_09460_),
    .Y(_09462_));
 sky130_fd_sc_hd__a211o_1 _16015_ (.A1(latched_is_lh),
    .A2(_09459_),
    .B1(_09462_),
    .C1(_09159_),
    .X(_09463_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16016_ (.A(_09463_),
    .X(_09464_));
 sky130_fd_sc_hd__o211a_1 _16017_ (.A1(_09459_),
    .A2(_09461_),
    .B1(_09464_),
    .C1(_08671_),
    .X(_09465_));
 sky130_fd_sc_hd__a211o_1 _16018_ (.A1(_08902_),
    .A2(_09457_),
    .B1(_09465_),
    .C1(_08666_),
    .X(_09466_));
 sky130_fd_sc_hd__o32a_1 _16019_ (.A1(_09429_),
    .A2(_09456_),
    .A3(_09466_),
    .B1(_09217_),
    .B2(\irq_pending[15] ),
    .X(_14578_));
 sky130_fd_sc_hd__or2_1 _16020_ (.A(\reg_pc[16] ),
    .B(\decoded_imm[16] ),
    .X(_09467_));
 sky130_fd_sc_hd__clkbuf_2 _16021_ (.A(\reg_pc[16] ),
    .X(_09468_));
 sky130_fd_sc_hd__nand2_1 _16022_ (.A(_09468_),
    .B(\decoded_imm[16] ),
    .Y(_09469_));
 sky130_fd_sc_hd__and2_1 _16023_ (.A(_09467_),
    .B(_09469_),
    .X(_09470_));
 sky130_fd_sc_hd__a21oi_1 _16024_ (.A1(_09387_),
    .A2(_09391_),
    .B1(_09425_),
    .Y(_09471_));
 sky130_fd_sc_hd__or2_1 _16025_ (.A(_09424_),
    .B(_09471_),
    .X(_09472_));
 sky130_fd_sc_hd__or2_1 _16026_ (.A(_09470_),
    .B(_09472_),
    .X(_09473_));
 sky130_fd_sc_hd__nand2_1 _16027_ (.A(_09470_),
    .B(_09472_),
    .Y(_09474_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16028_ (.A(_09464_),
    .X(_09475_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16029_ (.A(_08673_),
    .X(_09476_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16030_ (.A(_09460_),
    .X(_09477_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16031_ (.A(_09477_),
    .X(_09478_));
 sky130_fd_sc_hd__a21o_1 _16032_ (.A1(net40),
    .A2(_09476_),
    .B1(_09478_),
    .X(_09479_));
 sky130_fd_sc_hd__mux2_2 _16033_ (.A0(\genblk1.pcpi_mul.rd[16] ),
    .A1(\genblk1.pcpi_mul.rd[48] ),
    .S(_08769_),
    .X(_09480_));
 sky130_fd_sc_hd__a22o_1 _16034_ (.A1(\irq_pending[16] ),
    .A2(_08665_),
    .B1(_09480_),
    .B2(_08886_),
    .X(_09481_));
 sky130_fd_sc_hd__clkbuf_2 _16035_ (.A(_08656_),
    .X(_09482_));
 sky130_fd_sc_hd__clkbuf_2 _16036_ (.A(_08653_),
    .X(_09483_));
 sky130_fd_sc_hd__a22o_1 _16037_ (.A1(\count_instr[48] ),
    .A2(_08942_),
    .B1(_09286_),
    .B2(\count_cycle[48] ),
    .X(_09484_));
 sky130_fd_sc_hd__a221o_1 _16038_ (.A1(\count_instr[16] ),
    .A2(_09482_),
    .B1(\count_cycle[16] ),
    .B2(_09483_),
    .C1(_09484_),
    .X(_09485_));
 sky130_fd_sc_hd__mux2_1 _16039_ (.A0(\cpuregs[18][16] ),
    .A1(\cpuregs[19][16] ),
    .S(_08561_),
    .X(_09486_));
 sky130_fd_sc_hd__or2_1 _16040_ (.A(\cpuregs[16][16] ),
    .B(_09181_),
    .X(_09487_));
 sky130_fd_sc_hd__o211a_1 _16041_ (.A1(\cpuregs[17][16] ),
    .A2(_09112_),
    .B1(_08950_),
    .C1(_09487_),
    .X(_09488_));
 sky130_fd_sc_hd__a21oi_1 _16042_ (.A1(_08553_),
    .A2(_09486_),
    .B1(_09488_),
    .Y(_09489_));
 sky130_fd_sc_hd__mux2_1 _16043_ (.A0(\cpuregs[10][16] ),
    .A1(\cpuregs[11][16] ),
    .S(_09083_),
    .X(_09490_));
 sky130_fd_sc_hd__mux2_1 _16044_ (.A0(\cpuregs[8][16] ),
    .A1(\cpuregs[9][16] ),
    .S(_09186_),
    .X(_09491_));
 sky130_fd_sc_hd__mux2_1 _16045_ (.A0(_09490_),
    .A1(_09491_),
    .S(_08586_),
    .X(_09492_));
 sky130_fd_sc_hd__mux2_1 _16046_ (.A0(\cpuregs[12][16] ),
    .A1(\cpuregs[13][16] ),
    .S(_08618_),
    .X(_09493_));
 sky130_fd_sc_hd__mux2_1 _16047_ (.A0(\cpuregs[14][16] ),
    .A1(\cpuregs[15][16] ),
    .S(_08595_),
    .X(_09494_));
 sky130_fd_sc_hd__or2_1 _16048_ (.A(_08593_),
    .B(_09494_),
    .X(_09495_));
 sky130_fd_sc_hd__o211a_1 _16049_ (.A1(_09123_),
    .A2(_09493_),
    .B1(_09495_),
    .C1(_08600_),
    .X(_09496_));
 sky130_fd_sc_hd__a211o_1 _16050_ (.A1(_09117_),
    .A2(_09492_),
    .B1(_09496_),
    .C1(_08605_),
    .X(_09497_));
 sky130_fd_sc_hd__mux2_1 _16051_ (.A0(\cpuregs[2][16] ),
    .A1(\cpuregs[3][16] ),
    .S(_09134_),
    .X(_09498_));
 sky130_fd_sc_hd__mux2_1 _16052_ (.A0(\cpuregs[0][16] ),
    .A1(\cpuregs[1][16] ),
    .S(_09136_),
    .X(_09499_));
 sky130_fd_sc_hd__mux2_1 _16053_ (.A0(_09498_),
    .A1(_09499_),
    .S(_09080_),
    .X(_09500_));
 sky130_fd_sc_hd__mux2_1 _16054_ (.A0(\cpuregs[4][16] ),
    .A1(\cpuregs[5][16] ),
    .S(_09197_),
    .X(_09501_));
 sky130_fd_sc_hd__mux2_1 _16055_ (.A0(\cpuregs[6][16] ),
    .A1(\cpuregs[7][16] ),
    .S(_08842_),
    .X(_09502_));
 sky130_fd_sc_hd__or2_1 _16056_ (.A(_08735_),
    .B(_09502_),
    .X(_09503_));
 sky130_fd_sc_hd__o211a_1 _16057_ (.A1(_09139_),
    .A2(_09501_),
    .B1(_09503_),
    .C1(_08620_),
    .X(_09504_));
 sky130_fd_sc_hd__a211o_1 _16058_ (.A1(_08608_),
    .A2(_09500_),
    .B1(_09504_),
    .C1(_09202_),
    .X(_09505_));
 sky130_fd_sc_hd__a21oi_2 _16059_ (.A1(_09497_),
    .A2(_09505_),
    .B1(_09148_),
    .Y(_09506_));
 sky130_fd_sc_hd__a211o_4 _16060_ (.A1(_08545_),
    .A2(_09489_),
    .B1(_09506_),
    .C1(_09150_),
    .X(_09507_));
 sky130_fd_sc_hd__a221o_1 _16061_ (.A1(\irq_mask[16] ),
    .A2(_08936_),
    .B1(\timer[16] ),
    .B2(_08641_),
    .C1(_08646_),
    .X(_09508_));
 sky130_fd_sc_hd__o21bai_1 _16062_ (.A1(_09259_),
    .A2(_09507_),
    .B1_N(_09508_),
    .Y(_09509_));
 sky130_fd_sc_hd__o211a_1 _16063_ (.A1(_09337_),
    .A2(_09485_),
    .B1(_09509_),
    .C1(_08293_),
    .X(_09510_));
 sky130_fd_sc_hd__a311o_1 _16064_ (.A1(_08896_),
    .A2(_09475_),
    .A3(_09479_),
    .B1(_09481_),
    .C1(_09510_),
    .X(_09511_));
 sky130_fd_sc_hd__a31o_1 _16065_ (.A1(_09101_),
    .A2(_09473_),
    .A3(_09474_),
    .B1(_09511_),
    .X(_14579_));
 sky130_fd_sc_hd__or2_1 _16066_ (.A(\reg_pc[17] ),
    .B(\decoded_imm[17] ),
    .X(_09512_));
 sky130_fd_sc_hd__nand2_1 _16067_ (.A(\reg_pc[17] ),
    .B(\decoded_imm[17] ),
    .Y(_09513_));
 sky130_fd_sc_hd__and2_1 _16068_ (.A(_09512_),
    .B(_09513_),
    .X(_09514_));
 sky130_fd_sc_hd__o211ai_1 _16069_ (.A1(_09424_),
    .A2(_09471_),
    .B1(_09514_),
    .C1(_09470_),
    .Y(_09515_));
 sky130_fd_sc_hd__or2b_1 _16070_ (.A(_09469_),
    .B_N(_09514_),
    .X(_09516_));
 sky130_fd_sc_hd__nand2_1 _16071_ (.A(_09469_),
    .B(_09474_),
    .Y(_09517_));
 sky130_fd_sc_hd__o21a_1 _16072_ (.A1(_09514_),
    .A2(_09517_),
    .B1(_08872_),
    .X(_09518_));
 sky130_fd_sc_hd__and3_1 _16073_ (.A(_09515_),
    .B(_09516_),
    .C(_09518_),
    .X(_09519_));
 sky130_fd_sc_hd__buf_2 _16074_ (.A(_08771_),
    .X(_09520_));
 sky130_fd_sc_hd__mux2_2 _16075_ (.A0(\genblk1.pcpi_mul.rd[17] ),
    .A1(\genblk1.pcpi_mul.rd[49] ),
    .S(_08900_),
    .X(_09521_));
 sky130_fd_sc_hd__clkbuf_4 _16076_ (.A(_08673_),
    .X(_09522_));
 sky130_fd_sc_hd__a21o_1 _16077_ (.A1(net41),
    .A2(_09522_),
    .B1(_09477_),
    .X(_09523_));
 sky130_fd_sc_hd__mux2_1 _16078_ (.A0(\cpuregs[18][17] ),
    .A1(\cpuregs[19][17] ),
    .S(_08574_),
    .X(_09524_));
 sky130_fd_sc_hd__or2_1 _16079_ (.A(\cpuregs[16][17] ),
    .B(_08783_),
    .X(_09525_));
 sky130_fd_sc_hd__o211a_1 _16080_ (.A1(\cpuregs[17][17] ),
    .A2(_08827_),
    .B1(_08732_),
    .C1(_09525_),
    .X(_09526_));
 sky130_fd_sc_hd__a21oi_1 _16081_ (.A1(_08948_),
    .A2(_09524_),
    .B1(_09526_),
    .Y(_09527_));
 sky130_fd_sc_hd__mux2_1 _16082_ (.A0(\cpuregs[6][17] ),
    .A1(\cpuregs[7][17] ),
    .S(_08695_),
    .X(_09528_));
 sky130_fd_sc_hd__or2_1 _16083_ (.A(_08857_),
    .B(_09528_),
    .X(_09529_));
 sky130_fd_sc_hd__mux2_1 _16084_ (.A0(\cpuregs[4][17] ),
    .A1(\cpuregs[5][17] ),
    .S(_08572_),
    .X(_09530_));
 sky130_fd_sc_hd__o21a_1 _16085_ (.A1(_08713_),
    .A2(_09530_),
    .B1(_08973_),
    .X(_09531_));
 sky130_fd_sc_hd__mux2_1 _16086_ (.A0(\cpuregs[2][17] ),
    .A1(\cpuregs[3][17] ),
    .S(_08918_),
    .X(_09532_));
 sky130_fd_sc_hd__mux2_1 _16087_ (.A0(\cpuregs[0][17] ),
    .A1(\cpuregs[1][17] ),
    .S(_08918_),
    .X(_09533_));
 sky130_fd_sc_hd__mux2_1 _16088_ (.A0(_09532_),
    .A1(_09533_),
    .S(_08917_),
    .X(_09534_));
 sky130_fd_sc_hd__a221o_1 _16089_ (.A1(_09529_),
    .A2(_09531_),
    .B1(_09534_),
    .B2(_09026_),
    .C1(_08861_),
    .X(_09535_));
 sky130_fd_sc_hd__mux2_1 _16090_ (.A0(\cpuregs[8][17] ),
    .A1(\cpuregs[9][17] ),
    .S(_08695_),
    .X(_09536_));
 sky130_fd_sc_hd__mux2_1 _16091_ (.A0(\cpuregs[10][17] ),
    .A1(\cpuregs[11][17] ),
    .S(_08695_),
    .X(_09537_));
 sky130_fd_sc_hd__mux2_1 _16092_ (.A0(_09536_),
    .A1(_09537_),
    .S(_08550_),
    .X(_09538_));
 sky130_fd_sc_hd__mux2_1 _16093_ (.A0(\cpuregs[12][17] ),
    .A1(\cpuregs[13][17] ),
    .S(_08963_),
    .X(_09539_));
 sky130_fd_sc_hd__mux2_1 _16094_ (.A0(\cpuregs[14][17] ),
    .A1(\cpuregs[15][17] ),
    .S(_08609_),
    .X(_09540_));
 sky130_fd_sc_hd__or2_1 _16095_ (.A(_08585_),
    .B(_09540_),
    .X(_09541_));
 sky130_fd_sc_hd__o211a_1 _16096_ (.A1(_08713_),
    .A2(_09539_),
    .B1(_09541_),
    .C1(_08973_),
    .X(_09542_));
 sky130_fd_sc_hd__a211o_1 _16097_ (.A1(_09026_),
    .A2(_09538_),
    .B1(_09542_),
    .C1(_08975_),
    .X(_09543_));
 sky130_fd_sc_hd__a21oi_1 _16098_ (.A1(_09535_),
    .A2(_09543_),
    .B1(_08544_),
    .Y(_09544_));
 sky130_fd_sc_hd__a211o_4 _16099_ (.A1(_08932_),
    .A2(_09527_),
    .B1(_09544_),
    .C1(_08864_),
    .X(_09545_));
 sky130_fd_sc_hd__nor2_1 _16100_ (.A(_08688_),
    .B(_09545_),
    .Y(_09546_));
 sky130_fd_sc_hd__a221o_1 _16101_ (.A1(\irq_mask[17] ),
    .A2(_08936_),
    .B1(\timer[17] ),
    .B2(_08641_),
    .C1(_08645_),
    .X(_09547_));
 sky130_fd_sc_hd__a22o_1 _16102_ (.A1(\count_instr[49] ),
    .A2(_08657_),
    .B1(_08804_),
    .B2(\count_cycle[49] ),
    .X(_09548_));
 sky130_fd_sc_hd__a221o_1 _16103_ (.A1(\count_instr[17] ),
    .A2(_08656_),
    .B1(\count_cycle[17] ),
    .B2(_08653_),
    .C1(_09548_),
    .X(_09549_));
 sky130_fd_sc_hd__o22a_1 _16104_ (.A1(_09546_),
    .A2(_09547_),
    .B1(_09549_),
    .B2(_08649_),
    .X(_09550_));
 sky130_fd_sc_hd__a32o_1 _16105_ (.A1(_08880_),
    .A2(_09464_),
    .A3(_09523_),
    .B1(_09550_),
    .B2(_08945_),
    .X(_09551_));
 sky130_fd_sc_hd__a211o_1 _16106_ (.A1(_09520_),
    .A2(_09521_),
    .B1(_09551_),
    .C1(_08810_),
    .X(_09552_));
 sky130_fd_sc_hd__o22a_1 _16107_ (.A1(\irq_pending[17] ),
    .A2(_09217_),
    .B1(_09519_),
    .B2(_09552_),
    .X(_14580_));
 sky130_fd_sc_hd__clkbuf_2 _16108_ (.A(_08873_),
    .X(_09553_));
 sky130_fd_sc_hd__and3_1 _16109_ (.A(_09513_),
    .B(_09515_),
    .C(_09516_),
    .X(_09554_));
 sky130_fd_sc_hd__or2_1 _16110_ (.A(\reg_pc[18] ),
    .B(\decoded_imm[18] ),
    .X(_09555_));
 sky130_fd_sc_hd__nand2_1 _16111_ (.A(\reg_pc[18] ),
    .B(\decoded_imm[18] ),
    .Y(_09556_));
 sky130_fd_sc_hd__nand2_1 _16112_ (.A(_09555_),
    .B(_09556_),
    .Y(_09557_));
 sky130_fd_sc_hd__nand2_1 _16113_ (.A(_09554_),
    .B(_09557_),
    .Y(_09558_));
 sky130_fd_sc_hd__or2_1 _16114_ (.A(_09554_),
    .B(_09557_),
    .X(_09559_));
 sky130_fd_sc_hd__a21o_1 _16115_ (.A1(net42),
    .A2(_09476_),
    .B1(_09478_),
    .X(_09560_));
 sky130_fd_sc_hd__mux2_2 _16116_ (.A0(\genblk1.pcpi_mul.rd[18] ),
    .A1(\genblk1.pcpi_mul.rd[50] ),
    .S(_08769_),
    .X(_09561_));
 sky130_fd_sc_hd__a22o_1 _16117_ (.A1(\irq_pending[18] ),
    .A2(_08665_),
    .B1(_09561_),
    .B2(_08288_),
    .X(_09562_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16118_ (.A(_08804_),
    .X(_09563_));
 sky130_fd_sc_hd__a22o_1 _16119_ (.A1(\count_instr[50] ),
    .A2(_08942_),
    .B1(_09563_),
    .B2(\count_cycle[50] ),
    .X(_09564_));
 sky130_fd_sc_hd__a221o_1 _16120_ (.A1(\count_instr[18] ),
    .A2(_09482_),
    .B1(\count_cycle[18] ),
    .B2(_09483_),
    .C1(_09564_),
    .X(_09565_));
 sky130_fd_sc_hd__clkbuf_2 _16121_ (.A(_08688_),
    .X(_09566_));
 sky130_fd_sc_hd__mux2_1 _16122_ (.A0(\cpuregs[18][18] ),
    .A1(\cpuregs[19][18] ),
    .S(_08561_),
    .X(_09567_));
 sky130_fd_sc_hd__or2_1 _16123_ (.A(\cpuregs[16][18] ),
    .B(_09181_),
    .X(_09568_));
 sky130_fd_sc_hd__o211a_1 _16124_ (.A1(\cpuregs[17][18] ),
    .A2(_09112_),
    .B1(_08950_),
    .C1(_09568_),
    .X(_09569_));
 sky130_fd_sc_hd__a21oi_1 _16125_ (.A1(_08553_),
    .A2(_09567_),
    .B1(_09569_),
    .Y(_09570_));
 sky130_fd_sc_hd__mux2_1 _16126_ (.A0(\cpuregs[8][18] ),
    .A1(\cpuregs[9][18] ),
    .S(_09083_),
    .X(_09571_));
 sky130_fd_sc_hd__mux2_1 _16127_ (.A0(\cpuregs[10][18] ),
    .A1(\cpuregs[11][18] ),
    .S(_09186_),
    .X(_09572_));
 sky130_fd_sc_hd__mux2_1 _16128_ (.A0(_09571_),
    .A1(_09572_),
    .S(_08851_),
    .X(_09573_));
 sky130_fd_sc_hd__mux2_1 _16129_ (.A0(\cpuregs[12][18] ),
    .A1(\cpuregs[13][18] ),
    .S(_08618_),
    .X(_09574_));
 sky130_fd_sc_hd__mux2_1 _16130_ (.A0(\cpuregs[14][18] ),
    .A1(\cpuregs[15][18] ),
    .S(_09127_),
    .X(_09575_));
 sky130_fd_sc_hd__or2_1 _16131_ (.A(_09126_),
    .B(_09575_),
    .X(_09576_));
 sky130_fd_sc_hd__o211a_1 _16132_ (.A1(_09123_),
    .A2(_09574_),
    .B1(_09576_),
    .C1(_09130_),
    .X(_09577_));
 sky130_fd_sc_hd__a211o_1 _16133_ (.A1(_09117_),
    .A2(_09573_),
    .B1(_09577_),
    .C1(_08605_),
    .X(_09578_));
 sky130_fd_sc_hd__buf_2 _16134_ (.A(_09087_),
    .X(_09579_));
 sky130_fd_sc_hd__mux2_1 _16135_ (.A0(\cpuregs[6][18] ),
    .A1(\cpuregs[7][18] ),
    .S(_09134_),
    .X(_09580_));
 sky130_fd_sc_hd__mux2_1 _16136_ (.A0(\cpuregs[4][18] ),
    .A1(\cpuregs[5][18] ),
    .S(_09136_),
    .X(_09581_));
 sky130_fd_sc_hd__mux2_1 _16137_ (.A0(_09580_),
    .A1(_09581_),
    .S(_09080_),
    .X(_09582_));
 sky130_fd_sc_hd__mux2_1 _16138_ (.A0(\cpuregs[0][18] ),
    .A1(\cpuregs[1][18] ),
    .S(_09197_),
    .X(_09583_));
 sky130_fd_sc_hd__mux2_1 _16139_ (.A0(\cpuregs[2][18] ),
    .A1(\cpuregs[3][18] ),
    .S(_09143_),
    .X(_09584_));
 sky130_fd_sc_hd__or2_1 _16140_ (.A(_09142_),
    .B(_09584_),
    .X(_09585_));
 sky130_fd_sc_hd__o211a_1 _16141_ (.A1(_09139_),
    .A2(_09583_),
    .B1(_09585_),
    .C1(_08580_),
    .X(_09586_));
 sky130_fd_sc_hd__a211o_1 _16142_ (.A1(_09579_),
    .A2(_09582_),
    .B1(_09586_),
    .C1(_09202_),
    .X(_09587_));
 sky130_fd_sc_hd__a21oi_2 _16143_ (.A1(_09578_),
    .A2(_09587_),
    .B1(_09148_),
    .Y(_09588_));
 sky130_fd_sc_hd__a211o_4 _16144_ (.A1(_08545_),
    .A2(_09570_),
    .B1(_09588_),
    .C1(_09150_),
    .X(_09589_));
 sky130_fd_sc_hd__a221o_1 _16145_ (.A1(\irq_mask[18] ),
    .A2(_08936_),
    .B1(\timer[18] ),
    .B2(_08641_),
    .C1(_08646_),
    .X(_09590_));
 sky130_fd_sc_hd__o21bai_1 _16146_ (.A1(_09566_),
    .A2(_09589_),
    .B1_N(_09590_),
    .Y(_09591_));
 sky130_fd_sc_hd__o211a_1 _16147_ (.A1(_09337_),
    .A2(_09565_),
    .B1(_09591_),
    .C1(_08293_),
    .X(_09592_));
 sky130_fd_sc_hd__a311o_1 _16148_ (.A1(_08896_),
    .A2(_09475_),
    .A3(_09560_),
    .B1(_09562_),
    .C1(_09592_),
    .X(_09593_));
 sky130_fd_sc_hd__a31o_1 _16149_ (.A1(_09553_),
    .A2(_09558_),
    .A3(_09559_),
    .B1(_09593_),
    .X(_14581_));
 sky130_fd_sc_hd__or2_1 _16150_ (.A(\reg_pc[19] ),
    .B(\decoded_imm[19] ),
    .X(_09594_));
 sky130_fd_sc_hd__nand2_1 _16151_ (.A(\reg_pc[19] ),
    .B(\decoded_imm[19] ),
    .Y(_09595_));
 sky130_fd_sc_hd__nand2_1 _16152_ (.A(_09594_),
    .B(_09595_),
    .Y(_09596_));
 sky130_fd_sc_hd__and2_1 _16153_ (.A(_09556_),
    .B(_09559_),
    .X(_09597_));
 sky130_fd_sc_hd__nand2_1 _16154_ (.A(_09596_),
    .B(_09597_),
    .Y(_09598_));
 sky130_fd_sc_hd__o211a_1 _16155_ (.A1(_09596_),
    .A2(_09597_),
    .B1(_09598_),
    .C1(_08894_),
    .X(_09599_));
 sky130_fd_sc_hd__clkbuf_2 _16156_ (.A(_08886_),
    .X(_09600_));
 sky130_fd_sc_hd__mux2_1 _16157_ (.A0(\genblk1.pcpi_mul.rd[19] ),
    .A1(\genblk1.pcpi_mul.rd[51] ),
    .S(_08900_),
    .X(_09601_));
 sky130_fd_sc_hd__a21o_1 _16158_ (.A1(_09600_),
    .A2(_09601_),
    .B1(_08810_),
    .X(_09602_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16159_ (.A(_09463_),
    .X(_09603_));
 sky130_fd_sc_hd__a21o_1 _16160_ (.A1(net43),
    .A2(_09476_),
    .B1(_09461_),
    .X(_09604_));
 sky130_fd_sc_hd__mux2_1 _16161_ (.A0(\cpuregs[18][19] ),
    .A1(\cpuregs[19][19] ),
    .S(_08904_),
    .X(_09605_));
 sky130_fd_sc_hd__or2_1 _16162_ (.A(\cpuregs[16][19] ),
    .B(_08574_),
    .X(_09606_));
 sky130_fd_sc_hd__o211a_1 _16163_ (.A1(\cpuregs[17][19] ),
    .A2(_08565_),
    .B1(_08570_),
    .C1(_09606_),
    .X(_09607_));
 sky130_fd_sc_hd__a21oi_1 _16164_ (.A1(_08693_),
    .A2(_09605_),
    .B1(_09607_),
    .Y(_09608_));
 sky130_fd_sc_hd__mux2_1 _16165_ (.A0(\cpuregs[6][19] ),
    .A1(\cpuregs[7][19] ),
    .S(_08582_),
    .X(_09609_));
 sky130_fd_sc_hd__or2_1 _16166_ (.A(_08736_),
    .B(_09609_),
    .X(_09610_));
 sky130_fd_sc_hd__mux2_1 _16167_ (.A0(\cpuregs[4][19] ),
    .A1(\cpuregs[5][19] ),
    .S(_08590_),
    .X(_09611_));
 sky130_fd_sc_hd__o21a_1 _16168_ (.A1(_08589_),
    .A2(_09611_),
    .B1(_08620_),
    .X(_09612_));
 sky130_fd_sc_hd__mux2_1 _16169_ (.A0(\cpuregs[2][19] ),
    .A1(\cpuregs[3][19] ),
    .S(_08833_),
    .X(_09613_));
 sky130_fd_sc_hd__mux2_1 _16170_ (.A0(\cpuregs[0][19] ),
    .A1(\cpuregs[1][19] ),
    .S(_08835_),
    .X(_09614_));
 sky130_fd_sc_hd__mux2_1 _16171_ (.A0(_09613_),
    .A1(_09614_),
    .S(_08613_),
    .X(_09615_));
 sky130_fd_sc_hd__a221o_1 _16172_ (.A1(_09610_),
    .A2(_09612_),
    .B1(_09615_),
    .B2(_09075_),
    .C1(_09202_),
    .X(_09616_));
 sky130_fd_sc_hd__mux2_1 _16173_ (.A0(\cpuregs[14][19] ),
    .A1(\cpuregs[15][19] ),
    .S(_09118_),
    .X(_09617_));
 sky130_fd_sc_hd__mux2_1 _16174_ (.A0(\cpuregs[12][19] ),
    .A1(\cpuregs[13][19] ),
    .S(_09062_),
    .X(_09618_));
 sky130_fd_sc_hd__mux2_1 _16175_ (.A0(_09617_),
    .A1(_09618_),
    .S(_09121_),
    .X(_09619_));
 sky130_fd_sc_hd__mux2_1 _16176_ (.A0(\cpuregs[8][19] ),
    .A1(\cpuregs[9][19] ),
    .S(_09124_),
    .X(_09620_));
 sky130_fd_sc_hd__mux2_1 _16177_ (.A0(\cpuregs[10][19] ),
    .A1(\cpuregs[11][19] ),
    .S(_09069_),
    .X(_09621_));
 sky130_fd_sc_hd__or2_1 _16178_ (.A(_09068_),
    .B(_09621_),
    .X(_09622_));
 sky130_fd_sc_hd__o211a_1 _16179_ (.A1(_09065_),
    .A2(_09620_),
    .B1(_09622_),
    .C1(_08707_),
    .X(_09623_));
 sky130_fd_sc_hd__a211o_1 _16180_ (.A1(_09579_),
    .A2(_09619_),
    .B1(_09623_),
    .C1(_09073_),
    .X(_09624_));
 sky130_fd_sc_hd__a21oi_1 _16181_ (.A1(_09616_),
    .A2(_09624_),
    .B1(_08627_),
    .Y(_09625_));
 sky130_fd_sc_hd__a211o_4 _16182_ (.A1(_08903_),
    .A2(_09608_),
    .B1(_09625_),
    .C1(_08634_),
    .X(_09626_));
 sky130_fd_sc_hd__nor2_1 _16183_ (.A(_09566_),
    .B(_09626_),
    .Y(_09627_));
 sky130_fd_sc_hd__a221o_1 _16184_ (.A1(\irq_mask[19] ),
    .A2(_09206_),
    .B1(\timer[19] ),
    .B2(_09207_),
    .C1(_08939_),
    .X(_09628_));
 sky130_fd_sc_hd__a22o_1 _16185_ (.A1(\count_instr[51] ),
    .A2(_08801_),
    .B1(_09563_),
    .B2(\count_cycle[51] ),
    .X(_09629_));
 sky130_fd_sc_hd__a221o_1 _16186_ (.A1(\count_instr[19] ),
    .A2(_09482_),
    .B1(\count_cycle[19] ),
    .B2(_09483_),
    .C1(_09629_),
    .X(_09630_));
 sky130_fd_sc_hd__o22a_1 _16187_ (.A1(_09627_),
    .A2(_09628_),
    .B1(_09630_),
    .B2(_08650_),
    .X(_09631_));
 sky130_fd_sc_hd__a32o_1 _16188_ (.A1(_08896_),
    .A2(_09603_),
    .A3(_09604_),
    .B1(_09631_),
    .B2(_09210_),
    .X(_09632_));
 sky130_fd_sc_hd__o32a_1 _16189_ (.A1(_09599_),
    .A2(_09602_),
    .A3(_09632_),
    .B1(_09217_),
    .B2(\irq_pending[19] ),
    .X(_14582_));
 sky130_fd_sc_hd__or2_1 _16190_ (.A(\reg_pc[20] ),
    .B(\decoded_imm[20] ),
    .X(_09633_));
 sky130_fd_sc_hd__clkbuf_2 _16191_ (.A(\reg_pc[20] ),
    .X(_09634_));
 sky130_fd_sc_hd__nand2_1 _16192_ (.A(_09634_),
    .B(\decoded_imm[20] ),
    .Y(_09635_));
 sky130_fd_sc_hd__nand2_1 _16193_ (.A(_09633_),
    .B(_09635_),
    .Y(_09636_));
 sky130_fd_sc_hd__a311o_1 _16194_ (.A1(_09513_),
    .A2(_09515_),
    .A3(_09516_),
    .B1(_09557_),
    .C1(_09596_),
    .X(_09637_));
 sky130_fd_sc_hd__o211a_1 _16195_ (.A1(_09556_),
    .A2(_09596_),
    .B1(_09637_),
    .C1(_09595_),
    .X(_09638_));
 sky130_fd_sc_hd__nand2_1 _16196_ (.A(_09636_),
    .B(_09638_),
    .Y(_09639_));
 sky130_fd_sc_hd__or2_1 _16197_ (.A(_09636_),
    .B(_09638_),
    .X(_09640_));
 sky130_fd_sc_hd__a21o_1 _16198_ (.A1(net45),
    .A2(_09476_),
    .B1(_09478_),
    .X(_09641_));
 sky130_fd_sc_hd__mux2_2 _16199_ (.A0(\genblk1.pcpi_mul.rd[20] ),
    .A1(\genblk1.pcpi_mul.rd[52] ),
    .S(_08769_),
    .X(_09642_));
 sky130_fd_sc_hd__a22o_1 _16200_ (.A1(\irq_pending[20] ),
    .A2(_08665_),
    .B1(_09642_),
    .B2(_08288_),
    .X(_09643_));
 sky130_fd_sc_hd__a22o_1 _16201_ (.A1(\count_instr[52] ),
    .A2(_08942_),
    .B1(_09563_),
    .B2(\count_cycle[52] ),
    .X(_09644_));
 sky130_fd_sc_hd__a221o_1 _16202_ (.A1(\count_instr[20] ),
    .A2(_09482_),
    .B1(\count_cycle[20] ),
    .B2(_09483_),
    .C1(_09644_),
    .X(_09645_));
 sky130_fd_sc_hd__mux2_1 _16203_ (.A0(\cpuregs[18][20] ),
    .A1(\cpuregs[19][20] ),
    .S(_09110_),
    .X(_09646_));
 sky130_fd_sc_hd__or2_1 _16204_ (.A(\cpuregs[16][20] ),
    .B(_09056_),
    .X(_09647_));
 sky130_fd_sc_hd__o211a_1 _16205_ (.A1(\cpuregs[17][20] ),
    .A2(_09055_),
    .B1(_08950_),
    .C1(_09647_),
    .X(_09648_));
 sky130_fd_sc_hd__a21oi_1 _16206_ (.A1(_08553_),
    .A2(_09646_),
    .B1(_09648_),
    .Y(_09649_));
 sky130_fd_sc_hd__mux2_1 _16207_ (.A0(\cpuregs[6][20] ),
    .A1(\cpuregs[7][20] ),
    .S(_08610_),
    .X(_09650_));
 sky130_fd_sc_hd__or2_1 _16208_ (.A(_08736_),
    .B(_09650_),
    .X(_09651_));
 sky130_fd_sc_hd__mux2_1 _16209_ (.A0(\cpuregs[4][20] ),
    .A1(\cpuregs[5][20] ),
    .S(_08840_),
    .X(_09652_));
 sky130_fd_sc_hd__o21a_1 _16210_ (.A1(_08839_),
    .A2(_09652_),
    .B1(_08859_),
    .X(_09653_));
 sky130_fd_sc_hd__mux2_1 _16211_ (.A0(\cpuregs[2][20] ),
    .A1(\cpuregs[3][20] ),
    .S(_09078_),
    .X(_09654_));
 sky130_fd_sc_hd__mux2_1 _16212_ (.A0(\cpuregs[0][20] ),
    .A1(\cpuregs[1][20] ),
    .S(_09264_),
    .X(_09655_));
 sky130_fd_sc_hd__mux2_1 _16213_ (.A0(_09654_),
    .A1(_09655_),
    .S(_09018_),
    .X(_09656_));
 sky130_fd_sc_hd__a221o_1 _16214_ (.A1(_09651_),
    .A2(_09653_),
    .B1(_09656_),
    .B2(_08954_),
    .C1(_08617_),
    .X(_09657_));
 sky130_fd_sc_hd__mux2_1 _16215_ (.A0(\cpuregs[8][20] ),
    .A1(\cpuregs[9][20] ),
    .S(_09076_),
    .X(_09658_));
 sky130_fd_sc_hd__mux2_1 _16216_ (.A0(\cpuregs[10][20] ),
    .A1(\cpuregs[11][20] ),
    .S(_09076_),
    .X(_09659_));
 sky130_fd_sc_hd__mux2_1 _16217_ (.A0(_09658_),
    .A1(_09659_),
    .S(_08967_),
    .X(_09660_));
 sky130_fd_sc_hd__mux2_1 _16218_ (.A0(\cpuregs[12][20] ),
    .A1(\cpuregs[13][20] ),
    .S(_09140_),
    .X(_09661_));
 sky130_fd_sc_hd__mux2_1 _16219_ (.A0(\cpuregs[14][20] ),
    .A1(\cpuregs[15][20] ),
    .S(_09143_),
    .X(_09662_));
 sky130_fd_sc_hd__or2_1 _16220_ (.A(_09142_),
    .B(_09662_),
    .X(_09663_));
 sky130_fd_sc_hd__o211a_1 _16221_ (.A1(_09082_),
    .A2(_09661_),
    .B1(_09663_),
    .C1(_09087_),
    .X(_09664_));
 sky130_fd_sc_hd__a211o_1 _16222_ (.A1(_09075_),
    .A2(_09660_),
    .B1(_09664_),
    .C1(_08847_),
    .X(_09665_));
 sky130_fd_sc_hd__a21oi_2 _16223_ (.A1(_09657_),
    .A2(_09665_),
    .B1(_09090_),
    .Y(_09666_));
 sky130_fd_sc_hd__a211o_4 _16224_ (.A1(_09108_),
    .A2(_09649_),
    .B1(_09666_),
    .C1(_09092_),
    .X(_09667_));
 sky130_fd_sc_hd__a221o_1 _16225_ (.A1(\irq_mask[20] ),
    .A2(_08936_),
    .B1(\timer[20] ),
    .B2(_08641_),
    .C1(_08646_),
    .X(_09668_));
 sky130_fd_sc_hd__o21bai_1 _16226_ (.A1(_09566_),
    .A2(_09667_),
    .B1_N(_09668_),
    .Y(_09669_));
 sky130_fd_sc_hd__o211a_1 _16227_ (.A1(_09337_),
    .A2(_09645_),
    .B1(_09669_),
    .C1(_08293_),
    .X(_09670_));
 sky130_fd_sc_hd__a311o_1 _16228_ (.A1(_08896_),
    .A2(_09475_),
    .A3(_09641_),
    .B1(_09643_),
    .C1(_09670_),
    .X(_09671_));
 sky130_fd_sc_hd__a31o_1 _16229_ (.A1(_09553_),
    .A2(_09639_),
    .A3(_09640_),
    .B1(_09671_),
    .X(_14584_));
 sky130_fd_sc_hd__or2_1 _16230_ (.A(\reg_pc[21] ),
    .B(\decoded_imm[21] ),
    .X(_09672_));
 sky130_fd_sc_hd__nand2_1 _16231_ (.A(\reg_pc[21] ),
    .B(\decoded_imm[21] ),
    .Y(_09673_));
 sky130_fd_sc_hd__nand2_1 _16232_ (.A(_09672_),
    .B(_09673_),
    .Y(_09674_));
 sky130_fd_sc_hd__o21ai_1 _16233_ (.A1(_09636_),
    .A2(_09638_),
    .B1(_09635_),
    .Y(_09675_));
 sky130_vsdinv _16234_ (.A(_09675_),
    .Y(_09676_));
 sky130_fd_sc_hd__nand2_1 _16235_ (.A(_09674_),
    .B(_09676_),
    .Y(_09677_));
 sky130_fd_sc_hd__o211a_1 _16236_ (.A1(_09674_),
    .A2(_09676_),
    .B1(_09677_),
    .C1(_08872_),
    .X(_09678_));
 sky130_fd_sc_hd__mux2_1 _16237_ (.A0(\genblk1.pcpi_mul.rd[21] ),
    .A1(\genblk1.pcpi_mul.rd[53] ),
    .S(_08900_),
    .X(_09679_));
 sky130_fd_sc_hd__a21o_1 _16238_ (.A1(_09600_),
    .A2(_09679_),
    .B1(_08666_),
    .X(_09680_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16239_ (.A(_08673_),
    .X(_09681_));
 sky130_fd_sc_hd__a21o_1 _16240_ (.A1(net46),
    .A2(_09681_),
    .B1(_09461_),
    .X(_09682_));
 sky130_fd_sc_hd__mux2_1 _16241_ (.A0(\cpuregs[18][21] ),
    .A1(\cpuregs[19][21] ),
    .S(_08904_),
    .X(_09683_));
 sky130_fd_sc_hd__or2_1 _16242_ (.A(\cpuregs[16][21] ),
    .B(_08574_),
    .X(_09684_));
 sky130_fd_sc_hd__o211a_1 _16243_ (.A1(\cpuregs[17][21] ),
    .A2(_08565_),
    .B1(_08570_),
    .C1(_09684_),
    .X(_09685_));
 sky130_fd_sc_hd__a21oi_1 _16244_ (.A1(_08693_),
    .A2(_09683_),
    .B1(_09685_),
    .Y(_09686_));
 sky130_fd_sc_hd__mux2_1 _16245_ (.A0(\cpuregs[2][21] ),
    .A1(\cpuregs[3][21] ),
    .S(_08840_),
    .X(_09687_));
 sky130_fd_sc_hd__mux2_1 _16246_ (.A0(\cpuregs[0][21] ),
    .A1(\cpuregs[1][21] ),
    .S(_08840_),
    .X(_09688_));
 sky130_fd_sc_hd__mux2_1 _16247_ (.A0(_09687_),
    .A1(_09688_),
    .S(_08731_),
    .X(_09689_));
 sky130_fd_sc_hd__mux2_1 _16248_ (.A0(\cpuregs[4][21] ),
    .A1(\cpuregs[5][21] ),
    .S(_08590_),
    .X(_09690_));
 sky130_fd_sc_hd__mux2_1 _16249_ (.A0(\cpuregs[6][21] ),
    .A1(\cpuregs[7][21] ),
    .S(_08621_),
    .X(_09691_));
 sky130_fd_sc_hd__or2_1 _16250_ (.A(_08568_),
    .B(_09691_),
    .X(_09692_));
 sky130_fd_sc_hd__o211a_1 _16251_ (.A1(_08551_),
    .A2(_09690_),
    .B1(_09692_),
    .C1(_08600_),
    .X(_09693_));
 sky130_fd_sc_hd__a211o_1 _16252_ (.A1(_08581_),
    .A2(_09689_),
    .B1(_09693_),
    .C1(_08740_),
    .X(_09694_));
 sky130_fd_sc_hd__mux2_1 _16253_ (.A0(\cpuregs[14][21] ),
    .A1(\cpuregs[15][21] ),
    .S(_09186_),
    .X(_09695_));
 sky130_fd_sc_hd__mux2_1 _16254_ (.A0(\cpuregs[12][21] ),
    .A1(\cpuregs[13][21] ),
    .S(_09062_),
    .X(_09696_));
 sky130_fd_sc_hd__mux2_1 _16255_ (.A0(_09695_),
    .A1(_09696_),
    .S(_09121_),
    .X(_09697_));
 sky130_fd_sc_hd__mux2_1 _16256_ (.A0(\cpuregs[8][21] ),
    .A1(\cpuregs[9][21] ),
    .S(_09066_),
    .X(_09698_));
 sky130_fd_sc_hd__mux2_1 _16257_ (.A0(\cpuregs[10][21] ),
    .A1(\cpuregs[11][21] ),
    .S(_09069_),
    .X(_09699_));
 sky130_fd_sc_hd__or2_1 _16258_ (.A(_09068_),
    .B(_09699_),
    .X(_09700_));
 sky130_fd_sc_hd__o211a_1 _16259_ (.A1(_09065_),
    .A2(_09698_),
    .B1(_09700_),
    .C1(_08707_),
    .X(_09701_));
 sky130_fd_sc_hd__a211o_1 _16260_ (.A1(_09579_),
    .A2(_09697_),
    .B1(_09701_),
    .C1(_09073_),
    .X(_09702_));
 sky130_fd_sc_hd__a21oi_1 _16261_ (.A1(_09694_),
    .A2(_09702_),
    .B1(_08627_),
    .Y(_09703_));
 sky130_fd_sc_hd__a211o_4 _16262_ (.A1(_08903_),
    .A2(_09686_),
    .B1(_09703_),
    .C1(_08634_),
    .X(_09704_));
 sky130_fd_sc_hd__nor2_1 _16263_ (.A(_09566_),
    .B(_09704_),
    .Y(_09705_));
 sky130_fd_sc_hd__a221o_1 _16264_ (.A1(\irq_mask[21] ),
    .A2(_09206_),
    .B1(\timer[21] ),
    .B2(_09207_),
    .C1(_08939_),
    .X(_09706_));
 sky130_fd_sc_hd__a22o_1 _16265_ (.A1(\count_instr[53] ),
    .A2(_08801_),
    .B1(_09563_),
    .B2(\count_cycle[53] ),
    .X(_09707_));
 sky130_fd_sc_hd__a221o_1 _16266_ (.A1(\count_instr[21] ),
    .A2(_09482_),
    .B1(\count_cycle[21] ),
    .B2(_09483_),
    .C1(_09707_),
    .X(_09708_));
 sky130_fd_sc_hd__o22a_1 _16267_ (.A1(_09705_),
    .A2(_09706_),
    .B1(_09708_),
    .B2(_08650_),
    .X(_09709_));
 sky130_fd_sc_hd__a32o_1 _16268_ (.A1(_09048_),
    .A2(_09603_),
    .A3(_09682_),
    .B1(_09709_),
    .B2(_09210_),
    .X(_09710_));
 sky130_fd_sc_hd__o32a_1 _16269_ (.A1(_09678_),
    .A2(_09680_),
    .A3(_09710_),
    .B1(_08541_),
    .B2(\irq_pending[21] ),
    .X(_14585_));
 sky130_fd_sc_hd__or2_1 _16270_ (.A(\reg_pc[22] ),
    .B(\decoded_imm[22] ),
    .X(_09711_));
 sky130_fd_sc_hd__clkbuf_2 _16271_ (.A(\reg_pc[22] ),
    .X(_09712_));
 sky130_fd_sc_hd__nand2_1 _16272_ (.A(_09712_),
    .B(\decoded_imm[22] ),
    .Y(_09713_));
 sky130_fd_sc_hd__nand2_1 _16273_ (.A(_09711_),
    .B(_09713_),
    .Y(_09714_));
 sky130_fd_sc_hd__a21bo_1 _16274_ (.A1(_09672_),
    .A2(_09675_),
    .B1_N(_09673_),
    .X(_09715_));
 sky130_fd_sc_hd__xnor2_1 _16275_ (.A(_09714_),
    .B(_09715_),
    .Y(_09716_));
 sky130_fd_sc_hd__clkbuf_2 _16276_ (.A(_09522_),
    .X(_09717_));
 sky130_fd_sc_hd__a21o_1 _16277_ (.A1(net47),
    .A2(_09717_),
    .B1(_09478_),
    .X(_09718_));
 sky130_fd_sc_hd__mux2_2 _16278_ (.A0(\genblk1.pcpi_mul.rd[22] ),
    .A1(\genblk1.pcpi_mul.rd[54] ),
    .S(_08884_),
    .X(_09719_));
 sky130_fd_sc_hd__a22o_1 _16279_ (.A1(\irq_pending[22] ),
    .A2(_08773_),
    .B1(_09719_),
    .B2(_08771_),
    .X(_09720_));
 sky130_fd_sc_hd__a22o_1 _16280_ (.A1(\count_instr[54] ),
    .A2(_09375_),
    .B1(_09286_),
    .B2(\count_cycle[54] ),
    .X(_09721_));
 sky130_fd_sc_hd__a221o_1 _16281_ (.A1(\count_instr[22] ),
    .A2(_09285_),
    .B1(\count_cycle[22] ),
    .B2(_08654_),
    .C1(_09721_),
    .X(_09722_));
 sky130_fd_sc_hd__mux2_1 _16282_ (.A0(\cpuregs[16][22] ),
    .A1(\cpuregs[17][22] ),
    .S(_09110_),
    .X(_09723_));
 sky130_fd_sc_hd__or2_1 _16283_ (.A(\cpuregs[18][22] ),
    .B(_09056_),
    .X(_09724_));
 sky130_fd_sc_hd__o211a_1 _16284_ (.A1(\cpuregs[19][22] ),
    .A2(_09055_),
    .B1(_09113_),
    .C1(_09724_),
    .X(_09725_));
 sky130_fd_sc_hd__a21oi_1 _16285_ (.A1(_09109_),
    .A2(_09723_),
    .B1(_09725_),
    .Y(_09726_));
 sky130_fd_sc_hd__mux2_1 _16286_ (.A0(\cpuregs[10][22] ),
    .A1(\cpuregs[11][22] ),
    .S(_09060_),
    .X(_09727_));
 sky130_fd_sc_hd__mux2_1 _16287_ (.A0(\cpuregs[8][22] ),
    .A1(\cpuregs[9][22] ),
    .S(_09062_),
    .X(_09728_));
 sky130_fd_sc_hd__mux2_1 _16288_ (.A0(_09727_),
    .A1(_09728_),
    .S(_09121_),
    .X(_09729_));
 sky130_fd_sc_hd__mux2_1 _16289_ (.A0(\cpuregs[12][22] ),
    .A1(\cpuregs[13][22] ),
    .S(_09066_),
    .X(_09730_));
 sky130_fd_sc_hd__mux2_1 _16290_ (.A0(\cpuregs[14][22] ),
    .A1(\cpuregs[15][22] ),
    .S(_09069_),
    .X(_09731_));
 sky130_fd_sc_hd__or2_1 _16291_ (.A(_09068_),
    .B(_09731_),
    .X(_09732_));
 sky130_fd_sc_hd__o211a_1 _16292_ (.A1(_09065_),
    .A2(_09730_),
    .B1(_09732_),
    .C1(_09130_),
    .X(_09733_));
 sky130_fd_sc_hd__a211o_1 _16293_ (.A1(_08831_),
    .A2(_09729_),
    .B1(_09733_),
    .C1(_09073_),
    .X(_09734_));
 sky130_fd_sc_hd__mux2_1 _16294_ (.A0(\cpuregs[2][22] ),
    .A1(\cpuregs[3][22] ),
    .S(_09076_),
    .X(_09735_));
 sky130_fd_sc_hd__mux2_1 _16295_ (.A0(\cpuregs[0][22] ),
    .A1(\cpuregs[1][22] ),
    .S(_09078_),
    .X(_09736_));
 sky130_fd_sc_hd__mux2_1 _16296_ (.A0(_09735_),
    .A1(_09736_),
    .S(_09080_),
    .X(_09737_));
 sky130_fd_sc_hd__mux2_1 _16297_ (.A0(\cpuregs[4][22] ),
    .A1(\cpuregs[5][22] ),
    .S(_09140_),
    .X(_09738_));
 sky130_fd_sc_hd__mux2_1 _16298_ (.A0(\cpuregs[6][22] ),
    .A1(\cpuregs[7][22] ),
    .S(_08911_),
    .X(_09739_));
 sky130_fd_sc_hd__or2_1 _16299_ (.A(_09142_),
    .B(_09739_),
    .X(_09740_));
 sky130_fd_sc_hd__o211a_1 _16300_ (.A1(_09082_),
    .A2(_09738_),
    .B1(_09740_),
    .C1(_09087_),
    .X(_09741_));
 sky130_fd_sc_hd__a211o_1 _16301_ (.A1(_09075_),
    .A2(_09737_),
    .B1(_09741_),
    .C1(_08617_),
    .X(_09742_));
 sky130_fd_sc_hd__a21oi_2 _16302_ (.A1(_09734_),
    .A2(_09742_),
    .B1(_09090_),
    .Y(_09743_));
 sky130_fd_sc_hd__a211o_4 _16303_ (.A1(_09108_),
    .A2(_09726_),
    .B1(_09743_),
    .C1(_09092_),
    .X(_09744_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16304_ (.A(_08640_),
    .X(_09745_));
 sky130_fd_sc_hd__a221o_1 _16305_ (.A1(\irq_mask[22] ),
    .A2(_08637_),
    .B1(\timer[22] ),
    .B2(_09745_),
    .C1(_08646_),
    .X(_09746_));
 sky130_fd_sc_hd__o21bai_1 _16306_ (.A1(_09259_),
    .A2(_09744_),
    .B1_N(_09746_),
    .Y(_09747_));
 sky130_fd_sc_hd__o211a_1 _16307_ (.A1(_09378_),
    .A2(_09722_),
    .B1(_09747_),
    .C1(_09252_),
    .X(_09748_));
 sky130_fd_sc_hd__a311o_1 _16308_ (.A1(_08231_),
    .A2(_09475_),
    .A3(_09718_),
    .B1(_09720_),
    .C1(_09748_),
    .X(_09749_));
 sky130_fd_sc_hd__a21o_1 _16309_ (.A1(_09101_),
    .A2(_09716_),
    .B1(_09749_),
    .X(_14586_));
 sky130_fd_sc_hd__clkbuf_2 _16310_ (.A(\reg_pc[23] ),
    .X(_09750_));
 sky130_fd_sc_hd__buf_2 _16311_ (.A(\decoded_imm[23] ),
    .X(_09751_));
 sky130_fd_sc_hd__or2_1 _16312_ (.A(_09750_),
    .B(_09751_),
    .X(_09752_));
 sky130_fd_sc_hd__nand2_1 _16313_ (.A(_09750_),
    .B(_09751_),
    .Y(_09753_));
 sky130_fd_sc_hd__a21bo_1 _16314_ (.A1(_09711_),
    .A2(_09715_),
    .B1_N(_09713_),
    .X(_09754_));
 sky130_fd_sc_hd__a21oi_1 _16315_ (.A1(_09752_),
    .A2(_09753_),
    .B1(_09754_),
    .Y(_09755_));
 sky130_fd_sc_hd__a311oi_2 _16316_ (.A1(_09752_),
    .A2(_09753_),
    .A3(_09754_),
    .B1(_09755_),
    .C1(_09299_),
    .Y(_09756_));
 sky130_fd_sc_hd__mux2_1 _16317_ (.A0(\genblk1.pcpi_mul.rd[23] ),
    .A1(\genblk1.pcpi_mul.rd[55] ),
    .S(_08900_),
    .X(_09757_));
 sky130_fd_sc_hd__a21o_1 _16318_ (.A1(_09600_),
    .A2(_09757_),
    .B1(_08666_),
    .X(_09758_));
 sky130_fd_sc_hd__a21o_1 _16319_ (.A1(net48),
    .A2(_09681_),
    .B1(_09461_),
    .X(_09759_));
 sky130_fd_sc_hd__mux2_1 _16320_ (.A0(\cpuregs[18][23] ),
    .A1(\cpuregs[19][23] ),
    .S(_08904_),
    .X(_09760_));
 sky130_fd_sc_hd__or2_1 _16321_ (.A(\cpuregs[16][23] ),
    .B(_08629_),
    .X(_09761_));
 sky130_fd_sc_hd__o211a_1 _16322_ (.A1(\cpuregs[17][23] ),
    .A2(_08700_),
    .B1(_08701_),
    .C1(_09761_),
    .X(_09762_));
 sky130_fd_sc_hd__a21oi_1 _16323_ (.A1(_08693_),
    .A2(_09760_),
    .B1(_09762_),
    .Y(_09763_));
 sky130_fd_sc_hd__mux2_1 _16324_ (.A0(\cpuregs[8][23] ),
    .A1(\cpuregs[9][23] ),
    .S(_08718_),
    .X(_09764_));
 sky130_fd_sc_hd__mux2_1 _16325_ (.A0(\cpuregs[10][23] ),
    .A1(\cpuregs[11][23] ),
    .S(_08718_),
    .X(_09765_));
 sky130_fd_sc_hd__mux2_1 _16326_ (.A0(_09764_),
    .A1(_09765_),
    .S(_08851_),
    .X(_09766_));
 sky130_fd_sc_hd__mux2_1 _16327_ (.A0(\cpuregs[12][23] ),
    .A1(\cpuregs[13][23] ),
    .S(_08912_),
    .X(_09767_));
 sky130_fd_sc_hd__mux2_1 _16328_ (.A0(\cpuregs[14][23] ),
    .A1(\cpuregs[15][23] ),
    .S(_08621_),
    .X(_09768_));
 sky130_fd_sc_hd__or2_1 _16329_ (.A(_08568_),
    .B(_09768_),
    .X(_09769_));
 sky130_fd_sc_hd__o211a_1 _16330_ (.A1(_08551_),
    .A2(_09767_),
    .B1(_09769_),
    .C1(_08921_),
    .X(_09770_));
 sky130_fd_sc_hd__a211o_1 _16331_ (.A1(_08581_),
    .A2(_09766_),
    .B1(_09770_),
    .C1(_08726_),
    .X(_09771_));
 sky130_fd_sc_hd__mux2_1 _16332_ (.A0(\cpuregs[2][23] ),
    .A1(\cpuregs[3][23] ),
    .S(_08840_),
    .X(_09772_));
 sky130_fd_sc_hd__or2_1 _16333_ (.A(_08736_),
    .B(_09772_),
    .X(_09773_));
 sky130_fd_sc_hd__mux2_1 _16334_ (.A0(\cpuregs[0][23] ),
    .A1(\cpuregs[1][23] ),
    .S(_08590_),
    .X(_09774_));
 sky130_fd_sc_hd__o21a_1 _16335_ (.A1(_08551_),
    .A2(_09774_),
    .B1(_08580_),
    .X(_09775_));
 sky130_fd_sc_hd__mux2_1 _16336_ (.A0(\cpuregs[6][23] ),
    .A1(\cpuregs[7][23] ),
    .S(_09197_),
    .X(_09776_));
 sky130_fd_sc_hd__mux2_1 _16337_ (.A0(\cpuregs[4][23] ),
    .A1(\cpuregs[5][23] ),
    .S(_09140_),
    .X(_09777_));
 sky130_fd_sc_hd__mux2_1 _16338_ (.A0(_09776_),
    .A1(_09777_),
    .S(_08586_),
    .X(_09778_));
 sky130_fd_sc_hd__a221o_1 _16339_ (.A1(_09773_),
    .A2(_09775_),
    .B1(_09778_),
    .B2(_09579_),
    .C1(_09132_),
    .X(_09779_));
 sky130_fd_sc_hd__a21oi_2 _16340_ (.A1(_09771_),
    .A2(_09779_),
    .B1(_08932_),
    .Y(_09780_));
 sky130_fd_sc_hd__a211o_4 _16341_ (.A1(_08903_),
    .A2(_09763_),
    .B1(_09780_),
    .C1(_08743_),
    .X(_09781_));
 sky130_fd_sc_hd__nor2_1 _16342_ (.A(_09566_),
    .B(_09781_),
    .Y(_09782_));
 sky130_fd_sc_hd__a221o_1 _16343_ (.A1(\irq_mask[23] ),
    .A2(_09206_),
    .B1(\timer[23] ),
    .B2(_09207_),
    .C1(_08939_),
    .X(_09783_));
 sky130_fd_sc_hd__a22o_1 _16344_ (.A1(\count_instr[55] ),
    .A2(_08801_),
    .B1(_09563_),
    .B2(\count_cycle[55] ),
    .X(_09784_));
 sky130_fd_sc_hd__a221o_1 _16345_ (.A1(\count_instr[23] ),
    .A2(_08803_),
    .B1(\count_cycle[23] ),
    .B2(_08747_),
    .C1(_09784_),
    .X(_09785_));
 sky130_fd_sc_hd__o22a_1 _16346_ (.A1(_09782_),
    .A2(_09783_),
    .B1(_09785_),
    .B2(_08650_),
    .X(_09786_));
 sky130_fd_sc_hd__a32o_1 _16347_ (.A1(_09048_),
    .A2(_09603_),
    .A3(_09759_),
    .B1(_09786_),
    .B2(_08180_),
    .X(_09787_));
 sky130_fd_sc_hd__o32a_1 _16348_ (.A1(_09756_),
    .A2(_09758_),
    .A3(_09787_),
    .B1(_08541_),
    .B2(\irq_pending[23] ),
    .X(_14587_));
 sky130_fd_sc_hd__clkbuf_2 _16349_ (.A(\reg_pc[24] ),
    .X(_09788_));
 sky130_fd_sc_hd__nand2_1 _16350_ (.A(_09788_),
    .B(\decoded_imm[24] ),
    .Y(_09789_));
 sky130_fd_sc_hd__or2_1 _16351_ (.A(\reg_pc[24] ),
    .B(\decoded_imm[24] ),
    .X(_09790_));
 sky130_fd_sc_hd__nand2_1 _16352_ (.A(_09789_),
    .B(_09790_),
    .Y(_09791_));
 sky130_fd_sc_hd__and2_1 _16353_ (.A(_09750_),
    .B(_09751_),
    .X(_09792_));
 sky130_fd_sc_hd__a21o_1 _16354_ (.A1(_09752_),
    .A2(_09754_),
    .B1(_09792_),
    .X(_09793_));
 sky130_fd_sc_hd__xnor2_1 _16355_ (.A(_09791_),
    .B(_09793_),
    .Y(_09794_));
 sky130_fd_sc_hd__a21o_1 _16356_ (.A1(net49),
    .A2(_09717_),
    .B1(_09478_),
    .X(_09795_));
 sky130_fd_sc_hd__mux2_2 _16357_ (.A0(\genblk1.pcpi_mul.rd[24] ),
    .A1(\genblk1.pcpi_mul.rd[56] ),
    .S(_08884_),
    .X(_09796_));
 sky130_fd_sc_hd__a22o_1 _16358_ (.A1(\irq_pending[24] ),
    .A2(_08665_),
    .B1(_09796_),
    .B2(_08771_),
    .X(_09797_));
 sky130_fd_sc_hd__a22o_1 _16359_ (.A1(\count_instr[56] ),
    .A2(_09375_),
    .B1(_09286_),
    .B2(\count_cycle[56] ),
    .X(_09798_));
 sky130_fd_sc_hd__a221o_1 _16360_ (.A1(\count_instr[24] ),
    .A2(_09285_),
    .B1(\count_cycle[24] ),
    .B2(_08654_),
    .C1(_09798_),
    .X(_09799_));
 sky130_fd_sc_hd__mux2_1 _16361_ (.A0(\cpuregs[16][24] ),
    .A1(\cpuregs[17][24] ),
    .S(_09110_),
    .X(_09800_));
 sky130_fd_sc_hd__or2_1 _16362_ (.A(\cpuregs[18][24] ),
    .B(_09181_),
    .X(_09801_));
 sky130_fd_sc_hd__o211a_1 _16363_ (.A1(\cpuregs[19][24] ),
    .A2(_09112_),
    .B1(_09113_),
    .C1(_09801_),
    .X(_09802_));
 sky130_fd_sc_hd__a21oi_1 _16364_ (.A1(_09109_),
    .A2(_09800_),
    .B1(_09802_),
    .Y(_09803_));
 sky130_fd_sc_hd__mux2_1 _16365_ (.A0(\cpuregs[14][24] ),
    .A1(\cpuregs[15][24] ),
    .S(_09118_),
    .X(_09804_));
 sky130_fd_sc_hd__mux2_1 _16366_ (.A0(\cpuregs[12][24] ),
    .A1(\cpuregs[13][24] ),
    .S(_09186_),
    .X(_09805_));
 sky130_fd_sc_hd__mux2_1 _16367_ (.A0(_09804_),
    .A1(_09805_),
    .S(_08586_),
    .X(_09806_));
 sky130_fd_sc_hd__mux2_1 _16368_ (.A0(\cpuregs[8][24] ),
    .A1(\cpuregs[9][24] ),
    .S(_09124_),
    .X(_09807_));
 sky130_fd_sc_hd__mux2_1 _16369_ (.A0(\cpuregs[10][24] ),
    .A1(\cpuregs[11][24] ),
    .S(_09127_),
    .X(_09808_));
 sky130_fd_sc_hd__or2_1 _16370_ (.A(_09126_),
    .B(_09808_),
    .X(_09809_));
 sky130_fd_sc_hd__o211a_1 _16371_ (.A1(_09123_),
    .A2(_09807_),
    .B1(_09809_),
    .C1(_08707_),
    .X(_09810_));
 sky130_fd_sc_hd__a211o_1 _16372_ (.A1(_09579_),
    .A2(_09806_),
    .B1(_09810_),
    .C1(_08605_),
    .X(_09811_));
 sky130_fd_sc_hd__mux2_1 _16373_ (.A0(\cpuregs[2][24] ),
    .A1(\cpuregs[3][24] ),
    .S(_09264_),
    .X(_09812_));
 sky130_fd_sc_hd__or2_1 _16374_ (.A(_08731_),
    .B(_09812_),
    .X(_09813_));
 sky130_fd_sc_hd__mux2_1 _16375_ (.A0(\cpuregs[0][24] ),
    .A1(\cpuregs[1][24] ),
    .S(_08835_),
    .X(_09814_));
 sky130_fd_sc_hd__o21a_1 _16376_ (.A1(_08851_),
    .A2(_09814_),
    .B1(_08607_),
    .X(_09815_));
 sky130_fd_sc_hd__mux2_1 _16377_ (.A0(\cpuregs[6][24] ),
    .A1(\cpuregs[7][24] ),
    .S(_08559_),
    .X(_09816_));
 sky130_fd_sc_hd__mux2_1 _16378_ (.A0(\cpuregs[4][24] ),
    .A1(\cpuregs[5][24] ),
    .S(_08559_),
    .X(_09817_));
 sky130_fd_sc_hd__mux2_1 _16379_ (.A0(_09816_),
    .A1(_09817_),
    .S(_09018_),
    .X(_09818_));
 sky130_fd_sc_hd__a221o_1 _16380_ (.A1(_09813_),
    .A2(_09815_),
    .B1(_09818_),
    .B2(_08860_),
    .C1(_08617_),
    .X(_09819_));
 sky130_fd_sc_hd__a21oi_2 _16381_ (.A1(_09811_),
    .A2(_09819_),
    .B1(_09148_),
    .Y(_09820_));
 sky130_fd_sc_hd__a211o_4 _16382_ (.A1(_09108_),
    .A2(_09803_),
    .B1(_09820_),
    .C1(_09150_),
    .X(_09821_));
 sky130_fd_sc_hd__a221o_1 _16383_ (.A1(\irq_mask[24] ),
    .A2(_08637_),
    .B1(\timer[24] ),
    .B2(_09745_),
    .C1(_08646_),
    .X(_09822_));
 sky130_fd_sc_hd__o21bai_1 _16384_ (.A1(_09259_),
    .A2(_09821_),
    .B1_N(_09822_),
    .Y(_09823_));
 sky130_fd_sc_hd__o211a_1 _16385_ (.A1(_08650_),
    .A2(_09799_),
    .B1(_09823_),
    .C1(_08293_),
    .X(_09824_));
 sky130_fd_sc_hd__a311o_1 _16386_ (.A1(_08231_),
    .A2(_09475_),
    .A3(_09795_),
    .B1(_09797_),
    .C1(_09824_),
    .X(_09825_));
 sky130_fd_sc_hd__a21o_1 _16387_ (.A1(_09101_),
    .A2(_09794_),
    .B1(_09825_),
    .X(_14588_));
 sky130_fd_sc_hd__a21bo_1 _16388_ (.A1(_09790_),
    .A2(_09793_),
    .B1_N(_09789_),
    .X(_09826_));
 sky130_fd_sc_hd__or2_1 _16389_ (.A(\reg_pc[25] ),
    .B(\decoded_imm[25] ),
    .X(_09827_));
 sky130_fd_sc_hd__nand2_1 _16390_ (.A(\reg_pc[25] ),
    .B(\decoded_imm[25] ),
    .Y(_09828_));
 sky130_fd_sc_hd__nand3_1 _16391_ (.A(_09826_),
    .B(_09827_),
    .C(_09828_),
    .Y(_09829_));
 sky130_fd_sc_hd__a21o_1 _16392_ (.A1(_09827_),
    .A2(_09828_),
    .B1(_09826_),
    .X(_09830_));
 sky130_fd_sc_hd__a21o_1 _16393_ (.A1(net50),
    .A2(_09476_),
    .B1(_09461_),
    .X(_09831_));
 sky130_fd_sc_hd__mux2_2 _16394_ (.A0(\genblk1.pcpi_mul.rd[25] ),
    .A1(\genblk1.pcpi_mul.rd[57] ),
    .S(_08769_),
    .X(_09832_));
 sky130_fd_sc_hd__a22o_1 _16395_ (.A1(\irq_pending[25] ),
    .A2(_08665_),
    .B1(_09832_),
    .B2(_08288_),
    .X(_09833_));
 sky130_fd_sc_hd__mux2_1 _16396_ (.A0(\cpuregs[16][25] ),
    .A1(\cpuregs[17][25] ),
    .S(_09110_),
    .X(_09834_));
 sky130_fd_sc_hd__or2_1 _16397_ (.A(\cpuregs[18][25] ),
    .B(_09056_),
    .X(_09835_));
 sky130_fd_sc_hd__o211a_1 _16398_ (.A1(\cpuregs[19][25] ),
    .A2(_09055_),
    .B1(_09113_),
    .C1(_09835_),
    .X(_09836_));
 sky130_fd_sc_hd__a21oi_1 _16399_ (.A1(_09109_),
    .A2(_09834_),
    .B1(_09836_),
    .Y(_09837_));
 sky130_fd_sc_hd__mux2_1 _16400_ (.A0(\cpuregs[2][25] ),
    .A1(\cpuregs[3][25] ),
    .S(_09118_),
    .X(_09838_));
 sky130_fd_sc_hd__mux2_1 _16401_ (.A0(\cpuregs[0][25] ),
    .A1(\cpuregs[1][25] ),
    .S(_09060_),
    .X(_09839_));
 sky130_fd_sc_hd__mux2_1 _16402_ (.A0(_09838_),
    .A1(_09839_),
    .S(_09121_),
    .X(_09840_));
 sky130_fd_sc_hd__mux2_1 _16403_ (.A0(\cpuregs[4][25] ),
    .A1(\cpuregs[5][25] ),
    .S(_09124_),
    .X(_09841_));
 sky130_fd_sc_hd__mux2_1 _16404_ (.A0(\cpuregs[6][25] ),
    .A1(\cpuregs[7][25] ),
    .S(_09127_),
    .X(_09842_));
 sky130_fd_sc_hd__or2_1 _16405_ (.A(_09126_),
    .B(_09842_),
    .X(_09843_));
 sky130_fd_sc_hd__o211a_1 _16406_ (.A1(_09065_),
    .A2(_09841_),
    .B1(_09843_),
    .C1(_09130_),
    .X(_09844_));
 sky130_fd_sc_hd__a211o_1 _16407_ (.A1(_09117_),
    .A2(_09840_),
    .B1(_09844_),
    .C1(_09132_),
    .X(_09845_));
 sky130_fd_sc_hd__mux2_1 _16408_ (.A0(\cpuregs[8][25] ),
    .A1(\cpuregs[9][25] ),
    .S(_09134_),
    .X(_09846_));
 sky130_fd_sc_hd__mux2_1 _16409_ (.A0(\cpuregs[10][25] ),
    .A1(\cpuregs[11][25] ),
    .S(_09136_),
    .X(_09847_));
 sky130_fd_sc_hd__mux2_1 _16410_ (.A0(_09846_),
    .A1(_09847_),
    .S(_08967_),
    .X(_09848_));
 sky130_fd_sc_hd__mux2_1 _16411_ (.A0(\cpuregs[12][25] ),
    .A1(\cpuregs[13][25] ),
    .S(_09140_),
    .X(_09849_));
 sky130_fd_sc_hd__mux2_1 _16412_ (.A0(\cpuregs[14][25] ),
    .A1(\cpuregs[15][25] ),
    .S(_09143_),
    .X(_09850_));
 sky130_fd_sc_hd__or2_1 _16413_ (.A(_09142_),
    .B(_09850_),
    .X(_09851_));
 sky130_fd_sc_hd__o211a_1 _16414_ (.A1(_09082_),
    .A2(_09849_),
    .B1(_09851_),
    .C1(_08620_),
    .X(_09852_));
 sky130_fd_sc_hd__a211o_1 _16415_ (.A1(_08608_),
    .A2(_09848_),
    .B1(_09852_),
    .C1(_08847_),
    .X(_09853_));
 sky130_fd_sc_hd__a21oi_2 _16416_ (.A1(_09845_),
    .A2(_09853_),
    .B1(_09090_),
    .Y(_09854_));
 sky130_fd_sc_hd__a211o_4 _16417_ (.A1(_09108_),
    .A2(_09837_),
    .B1(_09854_),
    .C1(_09092_),
    .X(_09855_));
 sky130_fd_sc_hd__nor2_1 _16418_ (.A(_09566_),
    .B(_09855_),
    .Y(_09856_));
 sky130_fd_sc_hd__a221o_1 _16419_ (.A1(\irq_mask[25] ),
    .A2(_08937_),
    .B1(\timer[25] ),
    .B2(_08938_),
    .C1(_08939_),
    .X(_09857_));
 sky130_fd_sc_hd__a22o_1 _16420_ (.A1(\count_instr[57] ),
    .A2(_08942_),
    .B1(_09563_),
    .B2(\count_cycle[57] ),
    .X(_09858_));
 sky130_fd_sc_hd__a221o_1 _16421_ (.A1(\count_instr[25] ),
    .A2(_09482_),
    .B1(\count_cycle[25] ),
    .B2(_09483_),
    .C1(_09858_),
    .X(_09859_));
 sky130_fd_sc_hd__o221a_1 _16422_ (.A1(_09856_),
    .A2(_09857_),
    .B1(_09859_),
    .B2(_09337_),
    .C1(_08945_),
    .X(_09860_));
 sky130_fd_sc_hd__a311o_1 _16423_ (.A1(_08896_),
    .A2(_09603_),
    .A3(_09831_),
    .B1(_09833_),
    .C1(_09860_),
    .X(_09861_));
 sky130_fd_sc_hd__a31o_1 _16424_ (.A1(_09553_),
    .A2(_09829_),
    .A3(_09830_),
    .B1(_09861_),
    .X(_14589_));
 sky130_fd_sc_hd__or2_1 _16425_ (.A(\irq_pending[26] ),
    .B(_08540_),
    .X(_09862_));
 sky130_fd_sc_hd__a21o_1 _16426_ (.A1(net51),
    .A2(_09476_),
    .B1(_09478_),
    .X(_09863_));
 sky130_fd_sc_hd__mux2_2 _16427_ (.A0(\genblk1.pcpi_mul.rd[26] ),
    .A1(\genblk1.pcpi_mul.rd[58] ),
    .S(_08683_),
    .X(_09864_));
 sky130_fd_sc_hd__a22o_1 _16428_ (.A1(\count_instr[58] ),
    .A2(_08657_),
    .B1(_08804_),
    .B2(\count_cycle[58] ),
    .X(_09865_));
 sky130_fd_sc_hd__a221o_1 _16429_ (.A1(\count_instr[26] ),
    .A2(_08941_),
    .B1(\count_cycle[26] ),
    .B2(_08653_),
    .C1(_09865_),
    .X(_09866_));
 sky130_fd_sc_hd__mux2_1 _16430_ (.A0(\cpuregs[18][26] ),
    .A1(\cpuregs[19][26] ),
    .S(_09181_),
    .X(_09867_));
 sky130_fd_sc_hd__or2_1 _16431_ (.A(\cpuregs[16][26] ),
    .B(_08719_),
    .X(_09868_));
 sky130_fd_sc_hd__o211a_1 _16432_ (.A1(\cpuregs[17][26] ),
    .A2(_08564_),
    .B1(_08732_),
    .C1(_09868_),
    .X(_09869_));
 sky130_fd_sc_hd__a21oi_1 _16433_ (.A1(_08552_),
    .A2(_09867_),
    .B1(_09869_),
    .Y(_09870_));
 sky130_fd_sc_hd__mux2_1 _16434_ (.A0(\cpuregs[14][26] ),
    .A1(\cpuregs[15][26] ),
    .S(_08918_),
    .X(_09871_));
 sky130_fd_sc_hd__mux2_1 _16435_ (.A0(\cpuregs[12][26] ),
    .A1(\cpuregs[13][26] ),
    .S(_08717_),
    .X(_09872_));
 sky130_fd_sc_hd__mux2_1 _16436_ (.A0(_09871_),
    .A1(_09872_),
    .S(_08568_),
    .X(_09873_));
 sky130_fd_sc_hd__mux2_1 _16437_ (.A0(\cpuregs[8][26] ),
    .A1(\cpuregs[9][26] ),
    .S(_08695_),
    .X(_09874_));
 sky130_fd_sc_hd__mux2_1 _16438_ (.A0(\cpuregs[10][26] ),
    .A1(\cpuregs[11][26] ),
    .S(_08694_),
    .X(_09875_));
 sky130_fd_sc_hd__or2_1 _16439_ (.A(_08585_),
    .B(_09875_),
    .X(_09876_));
 sky130_fd_sc_hd__o211a_1 _16440_ (.A1(_08713_),
    .A2(_09874_),
    .B1(_09876_),
    .C1(_08706_),
    .X(_09877_));
 sky130_fd_sc_hd__a211o_1 _16441_ (.A1(_08921_),
    .A2(_09873_),
    .B1(_09877_),
    .C1(_08604_),
    .X(_09878_));
 sky130_fd_sc_hd__mux2_1 _16442_ (.A0(\cpuregs[2][26] ),
    .A1(\cpuregs[3][26] ),
    .S(_08717_),
    .X(_09879_));
 sky130_fd_sc_hd__mux2_1 _16443_ (.A0(\cpuregs[0][26] ),
    .A1(\cpuregs[1][26] ),
    .S(_08717_),
    .X(_09880_));
 sky130_fd_sc_hd__mux2_1 _16444_ (.A0(_09879_),
    .A1(_09880_),
    .S(_08568_),
    .X(_09881_));
 sky130_fd_sc_hd__mux2_1 _16445_ (.A0(\cpuregs[4][26] ),
    .A1(\cpuregs[5][26] ),
    .S(_08918_),
    .X(_09882_));
 sky130_fd_sc_hd__mux2_1 _16446_ (.A0(\cpuregs[6][26] ),
    .A1(\cpuregs[7][26] ),
    .S(_08694_),
    .X(_09883_));
 sky130_fd_sc_hd__or2_1 _16447_ (.A(_08585_),
    .B(_09883_),
    .X(_09884_));
 sky130_fd_sc_hd__o211a_1 _16448_ (.A1(_08713_),
    .A2(_09882_),
    .B1(_09884_),
    .C1(_08973_),
    .X(_09885_));
 sky130_fd_sc_hd__a211o_1 _16449_ (.A1(_09026_),
    .A2(_09881_),
    .B1(_09885_),
    .C1(_08616_),
    .X(_09886_));
 sky130_fd_sc_hd__a21oi_1 _16450_ (.A1(_09878_),
    .A2(_09886_),
    .B1(_08626_),
    .Y(_09887_));
 sky130_fd_sc_hd__a211o_4 _16451_ (.A1(_08691_),
    .A2(_09870_),
    .B1(_09887_),
    .C1(_08633_),
    .X(_09888_));
 sky130_fd_sc_hd__a221o_1 _16452_ (.A1(\irq_mask[26] ),
    .A2(instr_maskirq),
    .B1(\timer[26] ),
    .B2(_08640_),
    .C1(_08645_),
    .X(_09889_));
 sky130_fd_sc_hd__o21bai_1 _16453_ (.A1(_08688_),
    .A2(_09888_),
    .B1_N(_09889_),
    .Y(_09890_));
 sky130_fd_sc_hd__o211a_1 _16454_ (.A1(_08649_),
    .A2(_09866_),
    .B1(_09890_),
    .C1(_08179_),
    .X(_09891_));
 sky130_fd_sc_hd__a211o_1 _16455_ (.A1(_08886_),
    .A2(_09864_),
    .B1(_09891_),
    .C1(_08773_),
    .X(_09892_));
 sky130_fd_sc_hd__a31o_1 _16456_ (.A1(_08231_),
    .A2(_09475_),
    .A3(_09863_),
    .B1(_09892_),
    .X(_09893_));
 sky130_fd_sc_hd__clkbuf_2 _16457_ (.A(\reg_pc[26] ),
    .X(_09894_));
 sky130_fd_sc_hd__nand2_1 _16458_ (.A(_09894_),
    .B(\decoded_imm[26] ),
    .Y(_09895_));
 sky130_fd_sc_hd__or2_1 _16459_ (.A(_09894_),
    .B(\decoded_imm[26] ),
    .X(_09896_));
 sky130_fd_sc_hd__nand2_1 _16460_ (.A(_09895_),
    .B(_09896_),
    .Y(_09897_));
 sky130_fd_sc_hd__a21boi_1 _16461_ (.A1(_09826_),
    .A2(_09827_),
    .B1_N(_09828_),
    .Y(_09898_));
 sky130_fd_sc_hd__xor2_1 _16462_ (.A(_09897_),
    .B(_09898_),
    .X(_09899_));
 sky130_fd_sc_hd__a22o_1 _16463_ (.A1(_09862_),
    .A2(_09893_),
    .B1(_09899_),
    .B2(_09101_),
    .X(_14590_));
 sky130_fd_sc_hd__o21a_1 _16464_ (.A1(_09897_),
    .A2(_09898_),
    .B1(_09895_),
    .X(_09900_));
 sky130_fd_sc_hd__nor2_1 _16465_ (.A(\reg_pc[27] ),
    .B(\decoded_imm[27] ),
    .Y(_09901_));
 sky130_fd_sc_hd__clkbuf_2 _16466_ (.A(\reg_pc[27] ),
    .X(_09902_));
 sky130_fd_sc_hd__and2_1 _16467_ (.A(_09902_),
    .B(\decoded_imm[27] ),
    .X(_09903_));
 sky130_fd_sc_hd__or3_1 _16468_ (.A(_09900_),
    .B(_09901_),
    .C(_09903_),
    .X(_09904_));
 sky130_fd_sc_hd__o21ai_1 _16469_ (.A1(_09901_),
    .A2(_09903_),
    .B1(_09900_),
    .Y(_09905_));
 sky130_fd_sc_hd__a22o_1 _16470_ (.A1(\count_instr[59] ),
    .A2(_08658_),
    .B1(_08805_),
    .B2(\count_cycle[59] ),
    .X(_09906_));
 sky130_fd_sc_hd__a221o_1 _16471_ (.A1(\count_instr[27] ),
    .A2(_08749_),
    .B1(\count_cycle[27] ),
    .B2(_09037_),
    .C1(_09906_),
    .X(_09907_));
 sky130_fd_sc_hd__mux2_1 _16472_ (.A0(\cpuregs[18][27] ),
    .A1(\cpuregs[19][27] ),
    .S(_08629_),
    .X(_09908_));
 sky130_fd_sc_hd__or2_1 _16473_ (.A(\cpuregs[16][27] ),
    .B(_08783_),
    .X(_09909_));
 sky130_fd_sc_hd__o211a_1 _16474_ (.A1(\cpuregs[17][27] ),
    .A2(_08827_),
    .B1(_08732_),
    .C1(_09909_),
    .X(_09910_));
 sky130_fd_sc_hd__a21oi_1 _16475_ (.A1(_08948_),
    .A2(_09908_),
    .B1(_09910_),
    .Y(_09911_));
 sky130_fd_sc_hd__mux2_1 _16476_ (.A0(\cpuregs[10][27] ),
    .A1(\cpuregs[11][27] ),
    .S(_08572_),
    .X(_09912_));
 sky130_fd_sc_hd__mux2_1 _16477_ (.A0(\cpuregs[8][27] ),
    .A1(\cpuregs[9][27] ),
    .S(_08572_),
    .X(_09913_));
 sky130_fd_sc_hd__mux2_1 _16478_ (.A0(_09912_),
    .A1(_09913_),
    .S(_08857_),
    .X(_09914_));
 sky130_fd_sc_hd__mux2_1 _16479_ (.A0(\cpuregs[12][27] ),
    .A1(\cpuregs[13][27] ),
    .S(_08854_),
    .X(_09915_));
 sky130_fd_sc_hd__mux2_1 _16480_ (.A0(\cpuregs[14][27] ),
    .A1(\cpuregs[15][27] ),
    .S(_08571_),
    .X(_09916_));
 sky130_fd_sc_hd__or2_1 _16481_ (.A(_08969_),
    .B(_09916_),
    .X(_09917_));
 sky130_fd_sc_hd__o211a_1 _16482_ (.A1(_08837_),
    .A2(_09915_),
    .B1(_09917_),
    .C1(_08859_),
    .X(_09918_));
 sky130_fd_sc_hd__a211o_1 _16483_ (.A1(_08954_),
    .A2(_09914_),
    .B1(_09918_),
    .C1(_08975_),
    .X(_09919_));
 sky130_fd_sc_hd__mux2_1 _16484_ (.A0(\cpuregs[2][27] ),
    .A1(\cpuregs[3][27] ),
    .S(_08963_),
    .X(_09920_));
 sky130_fd_sc_hd__mux2_1 _16485_ (.A0(\cpuregs[0][27] ),
    .A1(\cpuregs[1][27] ),
    .S(_08963_),
    .X(_09921_));
 sky130_fd_sc_hd__mux2_1 _16486_ (.A0(_09920_),
    .A1(_09921_),
    .S(_08917_),
    .X(_09922_));
 sky130_fd_sc_hd__mux2_1 _16487_ (.A0(\cpuregs[4][27] ),
    .A1(\cpuregs[5][27] ),
    .S(_08709_),
    .X(_09923_));
 sky130_fd_sc_hd__mux2_1 _16488_ (.A0(\cpuregs[6][27] ),
    .A1(\cpuregs[7][27] ),
    .S(_08832_),
    .X(_09924_));
 sky130_fd_sc_hd__or2_1 _16489_ (.A(_08969_),
    .B(_09924_),
    .X(_09925_));
 sky130_fd_sc_hd__o211a_1 _16490_ (.A1(_08967_),
    .A2(_09923_),
    .B1(_09925_),
    .C1(_08973_),
    .X(_09926_));
 sky130_fd_sc_hd__a211o_1 _16491_ (.A1(_09026_),
    .A2(_09922_),
    .B1(_09926_),
    .C1(_08861_),
    .X(_09927_));
 sky130_fd_sc_hd__a21oi_1 _16492_ (.A1(_09919_),
    .A2(_09927_),
    .B1(_08691_),
    .Y(_09928_));
 sky130_fd_sc_hd__a211o_4 _16493_ (.A1(_08932_),
    .A2(_09911_),
    .B1(_09928_),
    .C1(_08864_),
    .X(_09929_));
 sky130_fd_sc_hd__a221o_1 _16494_ (.A1(\irq_mask[27] ),
    .A2(_08937_),
    .B1(\timer[27] ),
    .B2(_08938_),
    .C1(_09095_),
    .X(_09930_));
 sky130_fd_sc_hd__o21bai_1 _16495_ (.A1(_09009_),
    .A2(_09929_),
    .B1_N(_09930_),
    .Y(_09931_));
 sky130_fd_sc_hd__o211a_1 _16496_ (.A1(_09378_),
    .A2(_09907_),
    .B1(_09931_),
    .C1(_09252_),
    .X(_09932_));
 sky130_fd_sc_hd__a21o_1 _16497_ (.A1(net52),
    .A2(_09681_),
    .B1(_09477_),
    .X(_09933_));
 sky130_fd_sc_hd__mux2_2 _16498_ (.A0(\genblk1.pcpi_mul.rd[27] ),
    .A1(\genblk1.pcpi_mul.rd[59] ),
    .S(_08683_),
    .X(_09934_));
 sky130_fd_sc_hd__a21o_1 _16499_ (.A1(_08685_),
    .A2(_09934_),
    .B1(_08664_),
    .X(_09935_));
 sky130_fd_sc_hd__a31o_1 _16500_ (.A1(_09048_),
    .A2(_09603_),
    .A3(_09933_),
    .B1(_09935_),
    .X(_09936_));
 sky130_fd_sc_hd__o22a_1 _16501_ (.A1(\irq_pending[27] ),
    .A2(_09107_),
    .B1(_09932_),
    .B2(_09936_),
    .X(_09937_));
 sky130_fd_sc_hd__a31o_1 _16502_ (.A1(_09553_),
    .A2(_09904_),
    .A3(_09905_),
    .B1(_09937_),
    .X(_14591_));
 sky130_fd_sc_hd__nand2_2 _16503_ (.A(\reg_pc[28] ),
    .B(\decoded_imm[28] ),
    .Y(_09938_));
 sky130_fd_sc_hd__or2_1 _16504_ (.A(\reg_pc[28] ),
    .B(\decoded_imm[28] ),
    .X(_09939_));
 sky130_fd_sc_hd__nor2_1 _16505_ (.A(_09900_),
    .B(_09901_),
    .Y(_09940_));
 sky130_fd_sc_hd__a211o_1 _16506_ (.A1(_09938_),
    .A2(_09939_),
    .B1(_09940_),
    .C1(_09903_),
    .X(_09941_));
 sky130_fd_sc_hd__o211ai_2 _16507_ (.A1(_09903_),
    .A2(_09940_),
    .B1(_09939_),
    .C1(_09938_),
    .Y(_09942_));
 sky130_fd_sc_hd__a22o_1 _16508_ (.A1(\count_instr[60] ),
    .A2(_09375_),
    .B1(_08805_),
    .B2(\count_cycle[60] ),
    .X(_09943_));
 sky130_fd_sc_hd__a221o_1 _16509_ (.A1(\count_instr[28] ),
    .A2(_08749_),
    .B1(\count_cycle[28] ),
    .B2(_09037_),
    .C1(_09943_),
    .X(_09944_));
 sky130_fd_sc_hd__mux2_1 _16510_ (.A0(\cpuregs[16][28] ),
    .A1(\cpuregs[17][28] ),
    .S(_08561_),
    .X(_09945_));
 sky130_fd_sc_hd__or2_1 _16511_ (.A(\cpuregs[18][28] ),
    .B(_09181_),
    .X(_09946_));
 sky130_fd_sc_hd__o211a_1 _16512_ (.A1(\cpuregs[19][28] ),
    .A2(_08565_),
    .B1(_09113_),
    .C1(_09946_),
    .X(_09947_));
 sky130_fd_sc_hd__a21oi_1 _16513_ (.A1(_09109_),
    .A2(_09945_),
    .B1(_09947_),
    .Y(_09948_));
 sky130_fd_sc_hd__mux2_1 _16514_ (.A0(\cpuregs[2][28] ),
    .A1(\cpuregs[3][28] ),
    .S(_09197_),
    .X(_09949_));
 sky130_fd_sc_hd__mux2_1 _16515_ (.A0(\cpuregs[0][28] ),
    .A1(\cpuregs[1][28] ),
    .S(_09140_),
    .X(_09950_));
 sky130_fd_sc_hd__mux2_1 _16516_ (.A0(_09949_),
    .A1(_09950_),
    .S(_08586_),
    .X(_09951_));
 sky130_fd_sc_hd__mux2_1 _16517_ (.A0(\cpuregs[4][28] ),
    .A1(\cpuregs[5][28] ),
    .S(_08618_),
    .X(_09952_));
 sky130_fd_sc_hd__mux2_1 _16518_ (.A0(\cpuregs[6][28] ),
    .A1(\cpuregs[7][28] ),
    .S(_08595_),
    .X(_09953_));
 sky130_fd_sc_hd__or2_1 _16519_ (.A(_08593_),
    .B(_09953_),
    .X(_09954_));
 sky130_fd_sc_hd__o211a_1 _16520_ (.A1(_08589_),
    .A2(_09952_),
    .B1(_09954_),
    .C1(_08600_),
    .X(_09955_));
 sky130_fd_sc_hd__a211o_1 _16521_ (.A1(_08581_),
    .A2(_09951_),
    .B1(_09955_),
    .C1(_09132_),
    .X(_09956_));
 sky130_fd_sc_hd__mux2_1 _16522_ (.A0(\cpuregs[8][28] ),
    .A1(\cpuregs[9][28] ),
    .S(_08610_),
    .X(_09957_));
 sky130_fd_sc_hd__mux2_1 _16523_ (.A0(\cpuregs[10][28] ),
    .A1(\cpuregs[11][28] ),
    .S(_08610_),
    .X(_09958_));
 sky130_fd_sc_hd__mux2_1 _16524_ (.A0(_09957_),
    .A1(_09958_),
    .S(_08967_),
    .X(_09959_));
 sky130_fd_sc_hd__mux2_1 _16525_ (.A0(\cpuregs[12][28] ),
    .A1(\cpuregs[13][28] ),
    .S(_08582_),
    .X(_09960_));
 sky130_fd_sc_hd__mux2_1 _16526_ (.A0(\cpuregs[14][28] ),
    .A1(\cpuregs[15][28] ),
    .S(_08842_),
    .X(_09961_));
 sky130_fd_sc_hd__or2_1 _16527_ (.A(_08735_),
    .B(_09961_),
    .X(_09962_));
 sky130_fd_sc_hd__o211a_1 _16528_ (.A1(_09139_),
    .A2(_09960_),
    .B1(_09962_),
    .C1(_08620_),
    .X(_09963_));
 sky130_fd_sc_hd__a211o_1 _16529_ (.A1(_08608_),
    .A2(_09959_),
    .B1(_09963_),
    .C1(_08847_),
    .X(_09964_));
 sky130_fd_sc_hd__a21oi_2 _16530_ (.A1(_09956_),
    .A2(_09964_),
    .B1(_08627_),
    .Y(_09965_));
 sky130_fd_sc_hd__a211o_4 _16531_ (.A1(_08545_),
    .A2(_09948_),
    .B1(_09965_),
    .C1(_08634_),
    .X(_09966_));
 sky130_fd_sc_hd__a221o_1 _16532_ (.A1(\irq_mask[28] ),
    .A2(_08637_),
    .B1(\timer[28] ),
    .B2(_09745_),
    .C1(_09095_),
    .X(_09967_));
 sky130_fd_sc_hd__o21bai_1 _16533_ (.A1(_09009_),
    .A2(_09966_),
    .B1_N(_09967_),
    .Y(_09968_));
 sky130_fd_sc_hd__o211a_1 _16534_ (.A1(_09378_),
    .A2(_09944_),
    .B1(_09968_),
    .C1(_09252_),
    .X(_09969_));
 sky130_fd_sc_hd__a21o_1 _16535_ (.A1(net53),
    .A2(_09681_),
    .B1(_09477_),
    .X(_09970_));
 sky130_fd_sc_hd__mux2_2 _16536_ (.A0(\genblk1.pcpi_mul.rd[28] ),
    .A1(\genblk1.pcpi_mul.rd[60] ),
    .S(_08768_),
    .X(_09971_));
 sky130_fd_sc_hd__a21o_1 _16537_ (.A1(_08685_),
    .A2(_09971_),
    .B1(_08664_),
    .X(_09972_));
 sky130_fd_sc_hd__a31o_1 _16538_ (.A1(_08230_),
    .A2(_09464_),
    .A3(_09970_),
    .B1(_09972_),
    .X(_09973_));
 sky130_fd_sc_hd__o22a_1 _16539_ (.A1(\irq_pending[28] ),
    .A2(_09107_),
    .B1(_09969_),
    .B2(_09973_),
    .X(_09974_));
 sky130_fd_sc_hd__a31o_1 _16540_ (.A1(_09553_),
    .A2(_09941_),
    .A3(_09942_),
    .B1(_09974_),
    .X(_14592_));
 sky130_fd_sc_hd__clkbuf_2 _16541_ (.A(\reg_pc[29] ),
    .X(_09975_));
 sky130_fd_sc_hd__nor2_1 _16542_ (.A(_09975_),
    .B(\decoded_imm[29] ),
    .Y(_09976_));
 sky130_fd_sc_hd__and2_1 _16543_ (.A(_09975_),
    .B(\decoded_imm[29] ),
    .X(_09977_));
 sky130_fd_sc_hd__a211o_1 _16544_ (.A1(_09938_),
    .A2(_09942_),
    .B1(_09976_),
    .C1(_09977_),
    .X(_09978_));
 sky130_fd_sc_hd__o211ai_1 _16545_ (.A1(_09976_),
    .A2(_09977_),
    .B1(_09938_),
    .C1(_09942_),
    .Y(_09979_));
 sky130_fd_sc_hd__a22o_1 _16546_ (.A1(\count_instr[61] ),
    .A2(_09375_),
    .B1(_08805_),
    .B2(\count_cycle[61] ),
    .X(_09980_));
 sky130_fd_sc_hd__a221o_1 _16547_ (.A1(\count_instr[29] ),
    .A2(_09285_),
    .B1(\count_cycle[29] ),
    .B2(_09037_),
    .C1(_09980_),
    .X(_09981_));
 sky130_fd_sc_hd__mux2_1 _16548_ (.A0(\cpuregs[18][29] ),
    .A1(\cpuregs[19][29] ),
    .S(_08629_),
    .X(_09982_));
 sky130_fd_sc_hd__or2_1 _16549_ (.A(\cpuregs[16][29] ),
    .B(_08783_),
    .X(_09983_));
 sky130_fd_sc_hd__o211a_1 _16550_ (.A1(\cpuregs[17][29] ),
    .A2(_08827_),
    .B1(_08732_),
    .C1(_09983_),
    .X(_09984_));
 sky130_fd_sc_hd__a21oi_1 _16551_ (.A1(_08948_),
    .A2(_09982_),
    .B1(_09984_),
    .Y(_09985_));
 sky130_fd_sc_hd__mux2_1 _16552_ (.A0(\cpuregs[2][29] ),
    .A1(\cpuregs[3][29] ),
    .S(_08572_),
    .X(_09986_));
 sky130_fd_sc_hd__mux2_1 _16553_ (.A0(\cpuregs[0][29] ),
    .A1(\cpuregs[1][29] ),
    .S(_08572_),
    .X(_09987_));
 sky130_fd_sc_hd__mux2_1 _16554_ (.A0(_09986_),
    .A1(_09987_),
    .S(_08857_),
    .X(_09988_));
 sky130_fd_sc_hd__mux2_1 _16555_ (.A0(\cpuregs[4][29] ),
    .A1(\cpuregs[5][29] ),
    .S(_08854_),
    .X(_09989_));
 sky130_fd_sc_hd__mux2_1 _16556_ (.A0(\cpuregs[6][29] ),
    .A1(\cpuregs[7][29] ),
    .S(_08571_),
    .X(_09990_));
 sky130_fd_sc_hd__or2_1 _16557_ (.A(_08969_),
    .B(_09990_),
    .X(_09991_));
 sky130_fd_sc_hd__o211a_1 _16558_ (.A1(_08837_),
    .A2(_09989_),
    .B1(_09991_),
    .C1(_08859_),
    .X(_09992_));
 sky130_fd_sc_hd__a211o_1 _16559_ (.A1(_08954_),
    .A2(_09988_),
    .B1(_09992_),
    .C1(_08861_),
    .X(_09993_));
 sky130_fd_sc_hd__mux2_1 _16560_ (.A0(\cpuregs[8][29] ),
    .A1(\cpuregs[9][29] ),
    .S(_08963_),
    .X(_09994_));
 sky130_fd_sc_hd__mux2_1 _16561_ (.A0(\cpuregs[10][29] ),
    .A1(\cpuregs[11][29] ),
    .S(_08695_),
    .X(_09995_));
 sky130_fd_sc_hd__mux2_1 _16562_ (.A0(_09994_),
    .A1(_09995_),
    .S(_08550_),
    .X(_09996_));
 sky130_fd_sc_hd__mux2_1 _16563_ (.A0(\cpuregs[12][29] ),
    .A1(\cpuregs[13][29] ),
    .S(_08709_),
    .X(_09997_));
 sky130_fd_sc_hd__mux2_1 _16564_ (.A0(\cpuregs[14][29] ),
    .A1(\cpuregs[15][29] ),
    .S(_08832_),
    .X(_09998_));
 sky130_fd_sc_hd__or2_1 _16565_ (.A(_08969_),
    .B(_09998_),
    .X(_09999_));
 sky130_fd_sc_hd__o211a_1 _16566_ (.A1(_08713_),
    .A2(_09997_),
    .B1(_09999_),
    .C1(_08973_),
    .X(_10000_));
 sky130_fd_sc_hd__a211o_1 _16567_ (.A1(_09026_),
    .A2(_09996_),
    .B1(_10000_),
    .C1(_08975_),
    .X(_10001_));
 sky130_fd_sc_hd__a21oi_1 _16568_ (.A1(_09993_),
    .A2(_10001_),
    .B1(_08544_),
    .Y(_10002_));
 sky130_fd_sc_hd__a211o_4 _16569_ (.A1(_08932_),
    .A2(_09985_),
    .B1(_10002_),
    .C1(_08864_),
    .X(_10003_));
 sky130_fd_sc_hd__a221o_1 _16570_ (.A1(\irq_mask[29] ),
    .A2(_08637_),
    .B1(\timer[29] ),
    .B2(_09745_),
    .C1(_09095_),
    .X(_10004_));
 sky130_fd_sc_hd__o21bai_1 _16571_ (.A1(_09009_),
    .A2(_10003_),
    .B1_N(_10004_),
    .Y(_10005_));
 sky130_fd_sc_hd__o211a_1 _16572_ (.A1(_09378_),
    .A2(_09981_),
    .B1(_10005_),
    .C1(_09252_),
    .X(_10006_));
 sky130_fd_sc_hd__a21o_1 _16573_ (.A1(net54),
    .A2(_09681_),
    .B1(_09477_),
    .X(_10007_));
 sky130_fd_sc_hd__mux2_2 _16574_ (.A0(\genblk1.pcpi_mul.rd[29] ),
    .A1(\genblk1.pcpi_mul.rd[61] ),
    .S(_08768_),
    .X(_10008_));
 sky130_fd_sc_hd__a21o_1 _16575_ (.A1(_08685_),
    .A2(_10008_),
    .B1(_08664_),
    .X(_10009_));
 sky130_fd_sc_hd__a31o_1 _16576_ (.A1(_08230_),
    .A2(_09464_),
    .A3(_10007_),
    .B1(_10009_),
    .X(_10010_));
 sky130_fd_sc_hd__o22a_1 _16577_ (.A1(\irq_pending[29] ),
    .A2(_09107_),
    .B1(_10006_),
    .B2(_10010_),
    .X(_10011_));
 sky130_fd_sc_hd__a31o_1 _16578_ (.A1(_09553_),
    .A2(_09978_),
    .A3(_09979_),
    .B1(_10011_),
    .X(_14593_));
 sky130_fd_sc_hd__nand2_1 _16579_ (.A(\reg_pc[30] ),
    .B(\decoded_imm[30] ),
    .Y(_10012_));
 sky130_fd_sc_hd__or2_1 _16580_ (.A(\reg_pc[30] ),
    .B(\decoded_imm[30] ),
    .X(_10013_));
 sky130_fd_sc_hd__a21oi_1 _16581_ (.A1(_09938_),
    .A2(_09942_),
    .B1(_09976_),
    .Y(_10014_));
 sky130_fd_sc_hd__a211o_1 _16582_ (.A1(_10012_),
    .A2(_10013_),
    .B1(_10014_),
    .C1(_09977_),
    .X(_10015_));
 sky130_fd_sc_hd__o211ai_2 _16583_ (.A1(_09977_),
    .A2(_10014_),
    .B1(_10013_),
    .C1(_10012_),
    .Y(_10016_));
 sky130_fd_sc_hd__a22o_1 _16584_ (.A1(\count_instr[62] ),
    .A2(_09375_),
    .B1(_09286_),
    .B2(\count_cycle[62] ),
    .X(_10017_));
 sky130_fd_sc_hd__a221o_1 _16585_ (.A1(\count_instr[30] ),
    .A2(_09285_),
    .B1(\count_cycle[30] ),
    .B2(_08654_),
    .C1(_10017_),
    .X(_10018_));
 sky130_fd_sc_hd__mux2_1 _16586_ (.A0(\cpuregs[16][30] ),
    .A1(\cpuregs[17][30] ),
    .S(_09110_),
    .X(_10019_));
 sky130_fd_sc_hd__or2_1 _16587_ (.A(\cpuregs[18][30] ),
    .B(_09056_),
    .X(_10020_));
 sky130_fd_sc_hd__o211a_1 _16588_ (.A1(\cpuregs[19][30] ),
    .A2(_09112_),
    .B1(_09113_),
    .C1(_10020_),
    .X(_10021_));
 sky130_fd_sc_hd__a21oi_1 _16589_ (.A1(_09109_),
    .A2(_10019_),
    .B1(_10021_),
    .Y(_10022_));
 sky130_fd_sc_hd__mux2_1 _16590_ (.A0(\cpuregs[2][30] ),
    .A1(\cpuregs[3][30] ),
    .S(_09118_),
    .X(_10023_));
 sky130_fd_sc_hd__mux2_1 _16591_ (.A0(\cpuregs[0][30] ),
    .A1(\cpuregs[1][30] ),
    .S(_09186_),
    .X(_10024_));
 sky130_fd_sc_hd__mux2_1 _16592_ (.A0(_10023_),
    .A1(_10024_),
    .S(_09121_),
    .X(_10025_));
 sky130_fd_sc_hd__mux2_1 _16593_ (.A0(\cpuregs[4][30] ),
    .A1(\cpuregs[5][30] ),
    .S(_09124_),
    .X(_10026_));
 sky130_fd_sc_hd__mux2_1 _16594_ (.A0(\cpuregs[6][30] ),
    .A1(\cpuregs[7][30] ),
    .S(_09127_),
    .X(_10027_));
 sky130_fd_sc_hd__or2_1 _16595_ (.A(_09126_),
    .B(_10027_),
    .X(_10028_));
 sky130_fd_sc_hd__o211a_1 _16596_ (.A1(_09123_),
    .A2(_10026_),
    .B1(_10028_),
    .C1(_09130_),
    .X(_10029_));
 sky130_fd_sc_hd__a211o_1 _16597_ (.A1(_09117_),
    .A2(_10025_),
    .B1(_10029_),
    .C1(_09132_),
    .X(_10030_));
 sky130_fd_sc_hd__mux2_1 _16598_ (.A0(\cpuregs[14][30] ),
    .A1(\cpuregs[15][30] ),
    .S(_09134_),
    .X(_10031_));
 sky130_fd_sc_hd__mux2_1 _16599_ (.A0(\cpuregs[12][30] ),
    .A1(\cpuregs[13][30] ),
    .S(_09136_),
    .X(_10032_));
 sky130_fd_sc_hd__mux2_1 _16600_ (.A0(_10031_),
    .A1(_10032_),
    .S(_09080_),
    .X(_10033_));
 sky130_fd_sc_hd__mux2_1 _16601_ (.A0(\cpuregs[8][30] ),
    .A1(\cpuregs[9][30] ),
    .S(_09197_),
    .X(_10034_));
 sky130_fd_sc_hd__mux2_1 _16602_ (.A0(\cpuregs[10][30] ),
    .A1(\cpuregs[11][30] ),
    .S(_09143_),
    .X(_10035_));
 sky130_fd_sc_hd__or2_1 _16603_ (.A(_09142_),
    .B(_10035_),
    .X(_10036_));
 sky130_fd_sc_hd__o211a_1 _16604_ (.A1(_09139_),
    .A2(_10034_),
    .B1(_10036_),
    .C1(_08607_),
    .X(_10037_));
 sky130_fd_sc_hd__a211o_1 _16605_ (.A1(_09579_),
    .A2(_10033_),
    .B1(_10037_),
    .C1(_08847_),
    .X(_10038_));
 sky130_fd_sc_hd__a21oi_2 _16606_ (.A1(_10030_),
    .A2(_10038_),
    .B1(_09148_),
    .Y(_10039_));
 sky130_fd_sc_hd__a211o_4 _16607_ (.A1(_09108_),
    .A2(_10022_),
    .B1(_10039_),
    .C1(_09150_),
    .X(_10040_));
 sky130_fd_sc_hd__a221o_1 _16608_ (.A1(\irq_mask[30] ),
    .A2(_08637_),
    .B1(\timer[30] ),
    .B2(_09745_),
    .C1(_09095_),
    .X(_10041_));
 sky130_fd_sc_hd__o21bai_1 _16609_ (.A1(_09259_),
    .A2(_10040_),
    .B1_N(_10041_),
    .Y(_10042_));
 sky130_fd_sc_hd__o211a_1 _16610_ (.A1(_09378_),
    .A2(_10018_),
    .B1(_10042_),
    .C1(_09252_),
    .X(_10043_));
 sky130_fd_sc_hd__a21o_1 _16611_ (.A1(net56),
    .A2(_09522_),
    .B1(_09477_),
    .X(_10044_));
 sky130_fd_sc_hd__mux2_2 _16612_ (.A0(\genblk1.pcpi_mul.rd[30] ),
    .A1(\genblk1.pcpi_mul.rd[62] ),
    .S(_08768_),
    .X(_10045_));
 sky130_fd_sc_hd__a21o_1 _16613_ (.A1(_08287_),
    .A2(_10045_),
    .B1(_08664_),
    .X(_10046_));
 sky130_fd_sc_hd__a31o_1 _16614_ (.A1(_08230_),
    .A2(_09464_),
    .A3(_10044_),
    .B1(_10046_),
    .X(_10047_));
 sky130_fd_sc_hd__o22a_1 _16615_ (.A1(\irq_pending[30] ),
    .A2(_09107_),
    .B1(_10043_),
    .B2(_10047_),
    .X(_10048_));
 sky130_fd_sc_hd__a31o_1 _16616_ (.A1(_08873_),
    .A2(_10015_),
    .A3(_10016_),
    .B1(_10048_),
    .X(_14595_));
 sky130_fd_sc_hd__xnor2_1 _16617_ (.A(\reg_pc[31] ),
    .B(\decoded_imm[31] ),
    .Y(_10049_));
 sky130_fd_sc_hd__a21oi_1 _16618_ (.A1(_10012_),
    .A2(_10016_),
    .B1(_10049_),
    .Y(_10050_));
 sky130_fd_sc_hd__a31o_1 _16619_ (.A1(_10012_),
    .A2(_10016_),
    .A3(_10049_),
    .B1(_09299_),
    .X(_10051_));
 sky130_fd_sc_hd__a21o_1 _16620_ (.A1(net57),
    .A2(_09681_),
    .B1(_09461_),
    .X(_10052_));
 sky130_fd_sc_hd__mux2_2 _16621_ (.A0(\genblk1.pcpi_mul.rd[31] ),
    .A1(\genblk1.pcpi_mul.rd[63] ),
    .S(_08683_),
    .X(_10053_));
 sky130_fd_sc_hd__a22o_1 _16622_ (.A1(\count_instr[63] ),
    .A2(instr_rdinstrh),
    .B1(instr_rdcycleh),
    .B2(\count_cycle[63] ),
    .X(_10054_));
 sky130_fd_sc_hd__a221o_1 _16623_ (.A1(\count_instr[31] ),
    .A2(_08941_),
    .B1(\count_cycle[31] ),
    .B2(net373),
    .C1(_10054_),
    .X(_10055_));
 sky130_fd_sc_hd__mux2_1 _16624_ (.A0(\cpuregs[16][31] ),
    .A1(\cpuregs[17][31] ),
    .S(_08783_),
    .X(_10056_));
 sky130_fd_sc_hd__or2_1 _16625_ (.A(\cpuregs[18][31] ),
    .B(_08560_),
    .X(_10057_));
 sky130_fd_sc_hd__o211a_1 _16626_ (.A1(\cpuregs[19][31] ),
    .A2(_08564_),
    .B1(_08915_),
    .C1(_10057_),
    .X(_10058_));
 sky130_fd_sc_hd__a21oi_1 _16627_ (.A1(_08570_),
    .A2(_10056_),
    .B1(_10058_),
    .Y(_10059_));
 sky130_fd_sc_hd__mux2_1 _16628_ (.A0(\cpuregs[8][31] ),
    .A1(\cpuregs[9][31] ),
    .S(_08621_),
    .X(_10060_));
 sky130_fd_sc_hd__mux2_1 _16629_ (.A0(\cpuregs[10][31] ),
    .A1(\cpuregs[11][31] ),
    .S(_08621_),
    .X(_10061_));
 sky130_fd_sc_hd__mux2_1 _16630_ (.A0(_10060_),
    .A1(_10061_),
    .S(_08630_),
    .X(_10062_));
 sky130_fd_sc_hd__mux2_1 _16631_ (.A0(\cpuregs[12][31] ),
    .A1(\cpuregs[13][31] ),
    .S(_08621_),
    .X(_10063_));
 sky130_fd_sc_hd__mux2_1 _16632_ (.A0(\cpuregs[14][31] ),
    .A1(\cpuregs[15][31] ),
    .S(_08594_),
    .X(_10064_));
 sky130_fd_sc_hd__or2_1 _16633_ (.A(_08567_),
    .B(_10064_),
    .X(_10065_));
 sky130_fd_sc_hd__o211a_1 _16634_ (.A1(_08550_),
    .A2(_10063_),
    .B1(_10065_),
    .C1(_08599_),
    .X(_10066_));
 sky130_fd_sc_hd__a211o_1 _16635_ (.A1(_08707_),
    .A2(_10062_),
    .B1(_10066_),
    .C1(_08604_),
    .X(_10067_));
 sky130_fd_sc_hd__mux2_1 _16636_ (.A0(\cpuregs[0][31] ),
    .A1(\cpuregs[1][31] ),
    .S(_08842_),
    .X(_10068_));
 sky130_fd_sc_hd__or2_1 _16637_ (.A(_08588_),
    .B(_10068_),
    .X(_10069_));
 sky130_fd_sc_hd__mux2_1 _16638_ (.A0(\cpuregs[2][31] ),
    .A1(\cpuregs[3][31] ),
    .S(_08595_),
    .X(_10070_));
 sky130_fd_sc_hd__o21a_1 _16639_ (.A1(_08593_),
    .A2(_10070_),
    .B1(_08579_),
    .X(_10071_));
 sky130_fd_sc_hd__mux2_1 _16640_ (.A0(\cpuregs[6][31] ),
    .A1(\cpuregs[7][31] ),
    .S(_09143_),
    .X(_10072_));
 sky130_fd_sc_hd__mux2_1 _16641_ (.A0(\cpuregs[4][31] ),
    .A1(\cpuregs[5][31] ),
    .S(_08911_),
    .X(_10073_));
 sky130_fd_sc_hd__mux2_1 _16642_ (.A0(_10072_),
    .A1(_10073_),
    .S(_08730_),
    .X(_10074_));
 sky130_fd_sc_hd__a221o_1 _16643_ (.A1(_10069_),
    .A2(_10071_),
    .B1(_10074_),
    .B2(_09087_),
    .C1(_08616_),
    .X(_10075_));
 sky130_fd_sc_hd__a21oi_2 _16644_ (.A1(_10067_),
    .A2(_10075_),
    .B1(_08626_),
    .Y(_10076_));
 sky130_fd_sc_hd__a211o_4 _16645_ (.A1(_08544_),
    .A2(_10059_),
    .B1(_10076_),
    .C1(_08633_),
    .X(_10077_));
 sky130_fd_sc_hd__a221o_1 _16646_ (.A1(\irq_mask[31] ),
    .A2(instr_maskirq),
    .B1(\timer[31] ),
    .B2(_08640_),
    .C1(_08644_),
    .X(_10078_));
 sky130_fd_sc_hd__o21bai_1 _16647_ (.A1(_08688_),
    .A2(_10077_),
    .B1_N(_10078_),
    .Y(_10079_));
 sky130_fd_sc_hd__o211a_1 _16648_ (.A1(_08649_),
    .A2(_10055_),
    .B1(_10079_),
    .C1(_08178_),
    .X(_10080_));
 sky130_fd_sc_hd__a211o_1 _16649_ (.A1(_08685_),
    .A2(_10053_),
    .B1(_10080_),
    .C1(_08664_),
    .X(_10081_));
 sky130_fd_sc_hd__a31o_1 _16650_ (.A1(_09048_),
    .A2(_09603_),
    .A3(_10052_),
    .B1(_10081_),
    .X(_10082_));
 sky130_fd_sc_hd__o21ai_2 _16651_ (.A1(\irq_pending[31] ),
    .A2(_08541_),
    .B1(_10082_),
    .Y(_10083_));
 sky130_fd_sc_hd__o21ai_1 _16652_ (.A1(_10050_),
    .A2(_10051_),
    .B1(_10083_),
    .Y(_14596_));
 sky130_fd_sc_hd__or2_2 _16653_ (.A(instr_sll),
    .B(instr_slli),
    .X(_10084_));
 sky130_fd_sc_hd__or2_1 _16654_ (.A(instr_xor),
    .B(instr_xori),
    .X(_10085_));
 sky130_fd_sc_hd__or2_2 _16655_ (.A(instr_or),
    .B(instr_ori),
    .X(_10086_));
 sky130_fd_sc_hd__or2_2 _16656_ (.A(instr_and),
    .B(instr_andi),
    .X(_10087_));
 sky130_fd_sc_hd__or3_1 _16657_ (.A(_10085_),
    .B(_10086_),
    .C(_10087_),
    .X(_10088_));
 sky130_fd_sc_hd__or4_2 _16658_ (.A(is_compare),
    .B(_08218_),
    .C(_10084_),
    .D(_10088_),
    .X(_10089_));
 sky130_fd_sc_hd__buf_2 _16659_ (.A(_10089_),
    .X(_10090_));
 sky130_fd_sc_hd__buf_2 _16660_ (.A(_10090_),
    .X(_10091_));
 sky130_fd_sc_hd__nor4_1 _16661_ (.A(is_compare),
    .B(_08218_),
    .C(_10084_),
    .D(_10088_),
    .Y(_10092_));
 sky130_fd_sc_hd__clkbuf_2 _16662_ (.A(net371),
    .X(_10093_));
 sky130_fd_sc_hd__buf_2 _16663_ (.A(_10093_),
    .X(_10094_));
 sky130_fd_sc_hd__buf_2 _16664_ (.A(_08218_),
    .X(_10095_));
 sky130_fd_sc_hd__buf_2 _16665_ (.A(_10085_),
    .X(_10096_));
 sky130_fd_sc_hd__buf_2 _16666_ (.A(_10087_),
    .X(_10097_));
 sky130_fd_sc_hd__nor2_2 _16667_ (.A(instr_or),
    .B(instr_ori),
    .Y(_10098_));
 sky130_fd_sc_hd__nor2_1 _16668_ (.A(_08473_),
    .B(_10098_),
    .Y(_10099_));
 sky130_fd_sc_hd__a221o_1 _16669_ (.A1(\alu_shl[0] ),
    .A2(_10084_),
    .B1(_10097_),
    .B2(_08471_),
    .C1(_10099_),
    .X(_10100_));
 sky130_fd_sc_hd__a221o_1 _16670_ (.A1(\alu_shr[0] ),
    .A2(_10095_),
    .B1(_00000_),
    .B2(_10096_),
    .C1(_10100_),
    .X(_10101_));
 sky130_fd_sc_hd__a211o_1 _16671_ (.A1(is_compare),
    .A2(_08534_),
    .B1(_10094_),
    .C1(_10101_),
    .X(_10102_));
 sky130_fd_sc_hd__o21a_1 _16672_ (.A1(net429),
    .A2(_10091_),
    .B1(_10102_),
    .X(\alu_out[0] ));
 sky130_fd_sc_hd__clkbuf_2 _16673_ (.A(_10090_),
    .X(_10103_));
 sky130_fd_sc_hd__buf_4 _16674_ (.A(_08758_),
    .X(_10104_));
 sky130_fd_sc_hd__clkbuf_2 _16675_ (.A(net172),
    .X(_10105_));
 sky130_fd_sc_hd__clkbuf_2 _16676_ (.A(_10105_),
    .X(_10106_));
 sky130_fd_sc_hd__clkbuf_2 _16677_ (.A(_10106_),
    .X(_10107_));
 sky130_fd_sc_hd__clkbuf_8 _16678_ (.A(_10107_),
    .X(_10108_));
 sky130_fd_sc_hd__clkbuf_2 _16679_ (.A(_10087_),
    .X(_10109_));
 sky130_fd_sc_hd__buf_2 _16680_ (.A(_10109_),
    .X(_10110_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16681_ (.A(_10084_),
    .X(_10111_));
 sky130_fd_sc_hd__buf_2 _16682_ (.A(_10111_),
    .X(_10112_));
 sky130_fd_sc_hd__buf_2 _16683_ (.A(_10086_),
    .X(_10113_));
 sky130_fd_sc_hd__buf_2 _16684_ (.A(_10113_),
    .X(_10114_));
 sky130_fd_sc_hd__a22o_1 _16685_ (.A1(\alu_shl[1] ),
    .A2(_10112_),
    .B1(_10114_),
    .B2(_08465_),
    .X(_10115_));
 sky130_fd_sc_hd__a31o_1 _16686_ (.A1(_10104_),
    .A2(_10108_),
    .A3(_10110_),
    .B1(_10115_),
    .X(_10116_));
 sky130_fd_sc_hd__buf_2 _16687_ (.A(_08218_),
    .X(_10117_));
 sky130_fd_sc_hd__clkbuf_2 _16688_ (.A(_10117_),
    .X(_10118_));
 sky130_fd_sc_hd__buf_2 _16689_ (.A(_10096_),
    .X(_10119_));
 sky130_fd_sc_hd__clkbuf_2 _16690_ (.A(_10093_),
    .X(_10120_));
 sky130_fd_sc_hd__a221o_1 _16691_ (.A1(\alu_shr[1] ),
    .A2(_10118_),
    .B1(_08467_),
    .B2(_10119_),
    .C1(_10120_),
    .X(_10121_));
 sky130_fd_sc_hd__o22a_1 _16692_ (.A1(net431),
    .A2(_10103_),
    .B1(_10116_),
    .B2(_10121_),
    .X(\alu_out[1] ));
 sky130_fd_sc_hd__clkbuf_2 _16693_ (.A(_10111_),
    .X(_10122_));
 sky130_fd_sc_hd__buf_2 _16694_ (.A(_10109_),
    .X(_10123_));
 sky130_fd_sc_hd__and2_1 _16695_ (.A(net183),
    .B(_08456_),
    .X(_10124_));
 sky130_fd_sc_hd__a22o_1 _16696_ (.A1(_08454_),
    .A2(_10114_),
    .B1(_10123_),
    .B2(_10124_),
    .X(_10125_));
 sky130_fd_sc_hd__a21o_1 _16697_ (.A1(\alu_shl[2] ),
    .A2(_10122_),
    .B1(_10125_),
    .X(_10126_));
 sky130_fd_sc_hd__a221o_1 _16698_ (.A1(\alu_shr[2] ),
    .A2(_10118_),
    .B1(_08458_),
    .B2(_10119_),
    .C1(_10120_),
    .X(_10127_));
 sky130_fd_sc_hd__o22a_1 _16699_ (.A1(net426),
    .A2(_10103_),
    .B1(_10126_),
    .B2(_10127_),
    .X(\alu_out[2] ));
 sky130_fd_sc_hd__clkbuf_2 _16700_ (.A(_10111_),
    .X(_10128_));
 sky130_fd_sc_hd__buf_2 _16701_ (.A(_10085_),
    .X(_10129_));
 sky130_fd_sc_hd__and2_1 _16702_ (.A(net186),
    .B(net292),
    .X(_10130_));
 sky130_fd_sc_hd__a22o_1 _16703_ (.A1(_08442_),
    .A2(_10113_),
    .B1(_10097_),
    .B2(_10130_),
    .X(_10131_));
 sky130_fd_sc_hd__a221o_1 _16704_ (.A1(\alu_shl[3] ),
    .A2(_10128_),
    .B1(_10129_),
    .B2(_08445_),
    .C1(_10131_),
    .X(_10132_));
 sky130_fd_sc_hd__a211o_1 _16705_ (.A1(\alu_shr[3] ),
    .A2(_10118_),
    .B1(_10094_),
    .C1(_10132_),
    .X(_10133_));
 sky130_fd_sc_hd__o21a_1 _16706_ (.A1(net428),
    .A2(_10091_),
    .B1(_10133_),
    .X(\alu_out[3] ));
 sky130_fd_sc_hd__and2_1 _16707_ (.A(net187),
    .B(_08475_),
    .X(_10134_));
 sky130_fd_sc_hd__a22o_1 _16708_ (.A1(_08474_),
    .A2(_10114_),
    .B1(_10123_),
    .B2(_10134_),
    .X(_10135_));
 sky130_fd_sc_hd__a21o_1 _16709_ (.A1(\alu_shl[4] ),
    .A2(_10122_),
    .B1(_10135_),
    .X(_10136_));
 sky130_fd_sc_hd__a221o_1 _16710_ (.A1(\alu_shr[4] ),
    .A2(_10118_),
    .B1(_08477_),
    .B2(_10119_),
    .C1(_10120_),
    .X(_10137_));
 sky130_fd_sc_hd__o22a_1 _16711_ (.A1(net433),
    .A2(_10103_),
    .B1(_10136_),
    .B2(_10137_),
    .X(\alu_out[4] ));
 sky130_fd_sc_hd__a22o_1 _16712_ (.A1(_08450_),
    .A2(_10086_),
    .B1(_10097_),
    .B2(_08452_),
    .X(_10138_));
 sky130_fd_sc_hd__a221o_1 _16713_ (.A1(\alu_shr[5] ),
    .A2(_10095_),
    .B1(_10112_),
    .B2(\alu_shl[5] ),
    .C1(_10138_),
    .X(_10139_));
 sky130_fd_sc_hd__a211o_1 _16714_ (.A1(_08453_),
    .A2(_10119_),
    .B1(_10094_),
    .C1(_10139_),
    .X(_10140_));
 sky130_fd_sc_hd__o21a_1 _16715_ (.A1(net436),
    .A2(_10091_),
    .B1(_10140_),
    .X(\alu_out[5] ));
 sky130_fd_sc_hd__and2_1 _16716_ (.A(net189),
    .B(net295),
    .X(_10141_));
 sky130_fd_sc_hd__a22o_1 _16717_ (.A1(_08408_),
    .A2(_10086_),
    .B1(_10097_),
    .B2(_10141_),
    .X(_10142_));
 sky130_fd_sc_hd__a221o_1 _16718_ (.A1(\alu_shl[6] ),
    .A2(_10111_),
    .B1(_10096_),
    .B2(_08410_),
    .C1(_10142_),
    .X(_10143_));
 sky130_fd_sc_hd__a211o_1 _16719_ (.A1(\alu_shr[6] ),
    .A2(_10118_),
    .B1(_10094_),
    .C1(_10143_),
    .X(_10144_));
 sky130_fd_sc_hd__o21a_1 _16720_ (.A1(net442),
    .A2(_10091_),
    .B1(_10144_),
    .X(\alu_out[6] ));
 sky130_fd_sc_hd__or2_1 _16721_ (.A(net190),
    .B(net296),
    .X(_10145_));
 sky130_fd_sc_hd__a22o_1 _16722_ (.A1(_10145_),
    .A2(_10114_),
    .B1(_10123_),
    .B2(_08463_),
    .X(_10146_));
 sky130_fd_sc_hd__a21o_1 _16723_ (.A1(\alu_shl[7] ),
    .A2(_10122_),
    .B1(_10146_),
    .X(_10147_));
 sky130_fd_sc_hd__clkbuf_2 _16724_ (.A(_10096_),
    .X(_10148_));
 sky130_fd_sc_hd__a221o_1 _16725_ (.A1(\alu_shr[7] ),
    .A2(_10118_),
    .B1(_08464_),
    .B2(_10148_),
    .C1(_10120_),
    .X(_10149_));
 sky130_fd_sc_hd__o22a_1 _16726_ (.A1(net437),
    .A2(_10103_),
    .B1(_10147_),
    .B2(_10149_),
    .X(\alu_out[7] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16727_ (.A(_10098_),
    .X(_10150_));
 sky130_fd_sc_hd__buf_2 _16728_ (.A(_10150_),
    .X(_10151_));
 sky130_fd_sc_hd__a2bb2o_1 _16729_ (.A1_N(_08485_),
    .A2_N(_10151_),
    .B1(_10123_),
    .B2(_08483_),
    .X(_10152_));
 sky130_fd_sc_hd__a21o_1 _16730_ (.A1(\alu_shl[8] ),
    .A2(_10122_),
    .B1(_10152_),
    .X(_10153_));
 sky130_fd_sc_hd__clkbuf_2 _16731_ (.A(_10117_),
    .X(_10154_));
 sky130_fd_sc_hd__a221o_1 _16732_ (.A1(\alu_shr[8] ),
    .A2(_10154_),
    .B1(_08486_),
    .B2(_10148_),
    .C1(_10120_),
    .X(_10155_));
 sky130_fd_sc_hd__o22a_1 _16733_ (.A1(net430),
    .A2(_10103_),
    .B1(_10153_),
    .B2(_10155_),
    .X(\alu_out[8] ));
 sky130_fd_sc_hd__clkbuf_2 _16734_ (.A(net298),
    .X(_10156_));
 sky130_fd_sc_hd__clkbuf_4 _16735_ (.A(_10156_),
    .X(_10157_));
 sky130_fd_sc_hd__clkbuf_4 _16736_ (.A(net330),
    .X(_10158_));
 sky130_fd_sc_hd__a2bb2o_1 _16737_ (.A1_N(_08389_),
    .A2_N(_10151_),
    .B1(_10128_),
    .B2(\alu_shl[9] ),
    .X(_10159_));
 sky130_fd_sc_hd__a31o_1 _16738_ (.A1(_10157_),
    .A2(_10158_),
    .A3(_10110_),
    .B1(_10159_),
    .X(_10160_));
 sky130_fd_sc_hd__a221o_1 _16739_ (.A1(\alu_shr[9] ),
    .A2(_10154_),
    .B1(_08391_),
    .B2(_10148_),
    .C1(_10120_),
    .X(_10161_));
 sky130_fd_sc_hd__o22a_1 _16740_ (.A1(net434),
    .A2(_10103_),
    .B1(_10160_),
    .B2(_10161_),
    .X(\alu_out[9] ));
 sky130_fd_sc_hd__clkbuf_2 _16741_ (.A(_10090_),
    .X(_10162_));
 sky130_fd_sc_hd__clkbuf_4 _16742_ (.A(_08401_),
    .X(_10163_));
 sky130_fd_sc_hd__clkbuf_4 _16743_ (.A(net300),
    .X(_10164_));
 sky130_fd_sc_hd__buf_2 _16744_ (.A(_10111_),
    .X(_10165_));
 sky130_fd_sc_hd__a22o_1 _16745_ (.A1(\alu_shl[10] ),
    .A2(_10165_),
    .B1(_10114_),
    .B2(_08403_),
    .X(_10166_));
 sky130_fd_sc_hd__a31o_1 _16746_ (.A1(_10163_),
    .A2(_10164_),
    .A3(_10110_),
    .B1(_10166_),
    .X(_10167_));
 sky130_fd_sc_hd__clkbuf_2 _16747_ (.A(_10093_),
    .X(_10168_));
 sky130_fd_sc_hd__a221o_1 _16748_ (.A1(\alu_shr[10] ),
    .A2(_10154_),
    .B1(_08404_),
    .B2(_10148_),
    .C1(_10168_),
    .X(_10169_));
 sky130_fd_sc_hd__o22a_1 _16749_ (.A1(net445),
    .A2(_10162_),
    .B1(_10167_),
    .B2(_10169_),
    .X(\alu_out[10] ));
 sky130_fd_sc_hd__buf_2 _16750_ (.A(_10109_),
    .X(_10170_));
 sky130_fd_sc_hd__buf_2 _16751_ (.A(_10150_),
    .X(_10171_));
 sky130_fd_sc_hd__nor2_1 _16752_ (.A(_08415_),
    .B(_10171_),
    .Y(_10172_));
 sky130_fd_sc_hd__a221o_1 _16753_ (.A1(\alu_shl[11] ),
    .A2(_10122_),
    .B1(_10170_),
    .B2(_08414_),
    .C1(_10172_),
    .X(_10173_));
 sky130_fd_sc_hd__a221o_1 _16754_ (.A1(\alu_shr[11] ),
    .A2(_10154_),
    .B1(_08416_),
    .B2(_10148_),
    .C1(_10168_),
    .X(_10174_));
 sky130_fd_sc_hd__o22a_1 _16755_ (.A1(net435),
    .A2(_10162_),
    .B1(_10173_),
    .B2(_10174_),
    .X(\alu_out[11] ));
 sky130_fd_sc_hd__buf_2 _16756_ (.A(_10111_),
    .X(_10175_));
 sky130_fd_sc_hd__nor2_1 _16757_ (.A(_08344_),
    .B(_10171_),
    .Y(_10176_));
 sky130_fd_sc_hd__a221o_1 _16758_ (.A1(\alu_shl[12] ),
    .A2(_10175_),
    .B1(_10170_),
    .B2(_08341_),
    .C1(_10176_),
    .X(_10177_));
 sky130_fd_sc_hd__a221o_1 _16759_ (.A1(\alu_shr[12] ),
    .A2(_10154_),
    .B1(_08345_),
    .B2(_10148_),
    .C1(_10168_),
    .X(_10178_));
 sky130_fd_sc_hd__o22a_1 _16760_ (.A1(net432),
    .A2(_10162_),
    .B1(_10177_),
    .B2(_10178_),
    .X(\alu_out[12] ));
 sky130_fd_sc_hd__a2bb2o_1 _16761_ (.A1_N(_08348_),
    .A2_N(_10098_),
    .B1(_10097_),
    .B2(_08349_),
    .X(_10179_));
 sky130_fd_sc_hd__a221o_1 _16762_ (.A1(\alu_shr[13] ),
    .A2(_10117_),
    .B1(_10112_),
    .B2(\alu_shl[13] ),
    .C1(_10179_),
    .X(_10180_));
 sky130_fd_sc_hd__a211o_1 _16763_ (.A1(_08350_),
    .A2(_10119_),
    .B1(_10094_),
    .C1(_10180_),
    .X(_10181_));
 sky130_fd_sc_hd__o21a_1 _16764_ (.A1(net450),
    .A2(_10091_),
    .B1(_10181_),
    .X(\alu_out[13] ));
 sky130_fd_sc_hd__a2bb2o_1 _16765_ (.A1_N(_08420_),
    .A2_N(_10151_),
    .B1(_10109_),
    .B2(_08418_),
    .X(_10182_));
 sky130_fd_sc_hd__a21o_1 _16766_ (.A1(\alu_shl[14] ),
    .A2(_10122_),
    .B1(_10182_),
    .X(_10183_));
 sky130_fd_sc_hd__clkbuf_2 _16767_ (.A(_10096_),
    .X(_10184_));
 sky130_fd_sc_hd__a221o_1 _16768_ (.A1(\alu_shr[14] ),
    .A2(_10154_),
    .B1(_08421_),
    .B2(_10184_),
    .C1(_10168_),
    .X(_10185_));
 sky130_fd_sc_hd__o22a_1 _16769_ (.A1(net455),
    .A2(_10162_),
    .B1(_10183_),
    .B2(_10185_),
    .X(\alu_out[14] ));
 sky130_fd_sc_hd__clkbuf_2 _16770_ (.A(net273),
    .X(_10186_));
 sky130_fd_sc_hd__clkbuf_4 _16771_ (.A(_10186_),
    .X(_10187_));
 sky130_fd_sc_hd__clkbuf_4 _16772_ (.A(net305),
    .X(_10188_));
 sky130_fd_sc_hd__a2bb2o_1 _16773_ (.A1_N(_08446_),
    .A2_N(_10150_),
    .B1(_10128_),
    .B2(\alu_shl[15] ),
    .X(_10189_));
 sky130_fd_sc_hd__a31o_1 _16774_ (.A1(_10187_),
    .A2(_10188_),
    .A3(_10110_),
    .B1(_10189_),
    .X(_10190_));
 sky130_fd_sc_hd__clkbuf_2 _16775_ (.A(_10117_),
    .X(_10191_));
 sky130_fd_sc_hd__a221o_1 _16776_ (.A1(\alu_shr[15] ),
    .A2(_10191_),
    .B1(_08448_),
    .B2(_10184_),
    .C1(_10168_),
    .X(_10192_));
 sky130_fd_sc_hd__o22a_1 _16777_ (.A1(net465),
    .A2(_10162_),
    .B1(_10190_),
    .B2(_10192_),
    .X(\alu_out[15] ));
 sky130_fd_sc_hd__nor2_1 _16778_ (.A(_08380_),
    .B(_10171_),
    .Y(_10193_));
 sky130_fd_sc_hd__a221o_1 _16779_ (.A1(\alu_shl[16] ),
    .A2(_10175_),
    .B1(_10170_),
    .B2(_08379_),
    .C1(_10193_),
    .X(_10194_));
 sky130_fd_sc_hd__a221o_1 _16780_ (.A1(\alu_shr[16] ),
    .A2(_10191_),
    .B1(_08381_),
    .B2(_10184_),
    .C1(_10168_),
    .X(_10195_));
 sky130_fd_sc_hd__o22a_1 _16781_ (.A1(net427),
    .A2(_10162_),
    .B1(_10194_),
    .B2(_10195_),
    .X(\alu_out[16] ));
 sky130_fd_sc_hd__clkbuf_2 _16782_ (.A(_10090_),
    .X(_10196_));
 sky130_fd_sc_hd__clkbuf_4 _16783_ (.A(_08382_),
    .X(_10197_));
 sky130_fd_sc_hd__clkbuf_2 _16784_ (.A(_10109_),
    .X(_10198_));
 sky130_fd_sc_hd__a22o_1 _16785_ (.A1(\alu_shl[17] ),
    .A2(_10165_),
    .B1(_10114_),
    .B2(_08384_),
    .X(_10199_));
 sky130_fd_sc_hd__a31o_1 _16786_ (.A1(_10197_),
    .A2(_08383_),
    .A3(_10198_),
    .B1(_10199_),
    .X(_10200_));
 sky130_fd_sc_hd__clkbuf_2 _16787_ (.A(_10093_),
    .X(_10201_));
 sky130_fd_sc_hd__a221o_1 _16788_ (.A1(\alu_shr[17] ),
    .A2(_10191_),
    .B1(_08386_),
    .B2(_10184_),
    .C1(_10201_),
    .X(_10202_));
 sky130_fd_sc_hd__o22a_1 _16789_ (.A1(net425),
    .A2(_10196_),
    .B1(_10200_),
    .B2(_10202_),
    .X(\alu_out[17] ));
 sky130_fd_sc_hd__a2bb2o_1 _16790_ (.A1_N(_08353_),
    .A2_N(_10151_),
    .B1(_10175_),
    .B2(\alu_shl[18] ),
    .X(_10203_));
 sky130_fd_sc_hd__a21o_1 _16791_ (.A1(_08352_),
    .A2(_10110_),
    .B1(_10203_),
    .X(_10204_));
 sky130_fd_sc_hd__a221o_1 _16792_ (.A1(\alu_shr[18] ),
    .A2(_10191_),
    .B1(_08354_),
    .B2(_10184_),
    .C1(_10201_),
    .X(_10205_));
 sky130_fd_sc_hd__o22a_1 _16793_ (.A1(\alu_add_sub[18] ),
    .A2(_10196_),
    .B1(_10204_),
    .B2(_10205_),
    .X(\alu_out[18] ));
 sky130_fd_sc_hd__clkbuf_4 _16794_ (.A(_08374_),
    .X(_10206_));
 sky130_fd_sc_hd__a2bb2o_1 _16795_ (.A1_N(_08373_),
    .A2_N(_10150_),
    .B1(_10128_),
    .B2(\alu_shl[19] ),
    .X(_10207_));
 sky130_fd_sc_hd__a31o_1 _16796_ (.A1(_10206_),
    .A2(_08375_),
    .A3(_10198_),
    .B1(_10207_),
    .X(_10208_));
 sky130_fd_sc_hd__a221o_1 _16797_ (.A1(\alu_shr[19] ),
    .A2(_10191_),
    .B1(_08377_),
    .B2(_10184_),
    .C1(_10201_),
    .X(_10209_));
 sky130_fd_sc_hd__o22a_1 _16798_ (.A1(net460),
    .A2(_10196_),
    .B1(_10208_),
    .B2(_10209_),
    .X(\alu_out[19] ));
 sky130_fd_sc_hd__a2bb2o_1 _16799_ (.A1_N(_08357_),
    .A2_N(_10151_),
    .B1(_10112_),
    .B2(\alu_shl[20] ),
    .X(_10210_));
 sky130_fd_sc_hd__a21o_1 _16800_ (.A1(_08356_),
    .A2(_10110_),
    .B1(_10210_),
    .X(_10211_));
 sky130_fd_sc_hd__clkbuf_2 _16801_ (.A(_10096_),
    .X(_10212_));
 sky130_fd_sc_hd__a221o_1 _16802_ (.A1(\alu_shr[20] ),
    .A2(_10191_),
    .B1(_08358_),
    .B2(_10212_),
    .C1(_10201_),
    .X(_10213_));
 sky130_fd_sc_hd__o22a_1 _16803_ (.A1(net461),
    .A2(_10196_),
    .B1(_10211_),
    .B2(_10213_),
    .X(\alu_out[20] ));
 sky130_fd_sc_hd__buf_4 _16804_ (.A(_08363_),
    .X(_10214_));
 sky130_fd_sc_hd__a2bb2o_1 _16805_ (.A1_N(_08365_),
    .A2_N(_10150_),
    .B1(_10128_),
    .B2(\alu_shl[21] ),
    .X(_10215_));
 sky130_fd_sc_hd__a31o_1 _16806_ (.A1(_10214_),
    .A2(_08364_),
    .A3(_10198_),
    .B1(_10215_),
    .X(_10216_));
 sky130_fd_sc_hd__clkbuf_2 _16807_ (.A(_10117_),
    .X(_10217_));
 sky130_fd_sc_hd__a221o_1 _16808_ (.A1(\alu_shr[21] ),
    .A2(_10217_),
    .B1(_08367_),
    .B2(_10212_),
    .C1(_10201_),
    .X(_10218_));
 sky130_fd_sc_hd__o22a_1 _16809_ (.A1(\alu_add_sub[21] ),
    .A2(_10196_),
    .B1(_10216_),
    .B2(_10218_),
    .X(\alu_out[21] ));
 sky130_fd_sc_hd__nor2_1 _16810_ (.A(_08361_),
    .B(_10171_),
    .Y(_10219_));
 sky130_fd_sc_hd__a221o_1 _16811_ (.A1(\alu_shl[22] ),
    .A2(_10175_),
    .B1(_10170_),
    .B2(_08360_),
    .C1(_10219_),
    .X(_10220_));
 sky130_fd_sc_hd__a221o_1 _16812_ (.A1(\alu_shr[22] ),
    .A2(_10217_),
    .B1(_08362_),
    .B2(_10212_),
    .C1(_10201_),
    .X(_10221_));
 sky130_fd_sc_hd__o22a_1 _16813_ (.A1(net443),
    .A2(_10196_),
    .B1(_10220_),
    .B2(_10221_),
    .X(\alu_out[22] ));
 sky130_fd_sc_hd__clkbuf_2 _16814_ (.A(_10089_),
    .X(_10222_));
 sky130_fd_sc_hd__clkbuf_2 _16815_ (.A(net282),
    .X(_10223_));
 sky130_fd_sc_hd__clkbuf_4 _16816_ (.A(_10223_),
    .X(_10224_));
 sky130_fd_sc_hd__a32o_1 _16817_ (.A1(_10224_),
    .A2(_08369_),
    .A3(_10109_),
    .B1(_10112_),
    .B2(\alu_shl[23] ),
    .X(_10225_));
 sky130_fd_sc_hd__o21bai_1 _16818_ (.A1(_08368_),
    .A2(_10171_),
    .B1_N(_10225_),
    .Y(_10226_));
 sky130_fd_sc_hd__clkbuf_2 _16819_ (.A(net371),
    .X(_10227_));
 sky130_fd_sc_hd__a221o_1 _16820_ (.A1(\alu_shr[23] ),
    .A2(_10217_),
    .B1(_08371_),
    .B2(_10212_),
    .C1(_10227_),
    .X(_10228_));
 sky130_fd_sc_hd__o22a_1 _16821_ (.A1(\alu_add_sub[23] ),
    .A2(_10222_),
    .B1(_10226_),
    .B2(_10228_),
    .X(\alu_out[23] ));
 sky130_fd_sc_hd__nor2_1 _16822_ (.A(_08425_),
    .B(_10171_),
    .Y(_10229_));
 sky130_fd_sc_hd__a221o_1 _16823_ (.A1(\alu_shl[24] ),
    .A2(_10175_),
    .B1(_10123_),
    .B2(_08424_),
    .C1(_10229_),
    .X(_10230_));
 sky130_fd_sc_hd__a221o_1 _16824_ (.A1(\alu_shr[24] ),
    .A2(_10217_),
    .B1(_08426_),
    .B2(_10212_),
    .C1(_10227_),
    .X(_10231_));
 sky130_fd_sc_hd__o22a_1 _16825_ (.A1(net421),
    .A2(_10222_),
    .B1(_10230_),
    .B2(_10231_),
    .X(\alu_out[24] ));
 sky130_fd_sc_hd__clkbuf_2 _16826_ (.A(net284),
    .X(_10232_));
 sky130_fd_sc_hd__or2_1 _16827_ (.A(_10232_),
    .B(_08427_),
    .X(_10233_));
 sky130_fd_sc_hd__a22o_1 _16828_ (.A1(_10233_),
    .A2(_10086_),
    .B1(_10097_),
    .B2(_08429_),
    .X(_10234_));
 sky130_fd_sc_hd__a221o_1 _16829_ (.A1(\alu_shr[25] ),
    .A2(_10117_),
    .B1(_10112_),
    .B2(\alu_shl[25] ),
    .C1(_10234_),
    .X(_10235_));
 sky130_fd_sc_hd__a211o_1 _16830_ (.A1(_08430_),
    .A2(_10119_),
    .B1(_10094_),
    .C1(_10235_),
    .X(_10236_));
 sky130_fd_sc_hd__o21a_1 _16831_ (.A1(net424),
    .A2(_10091_),
    .B1(_10236_),
    .X(\alu_out[25] ));
 sky130_fd_sc_hd__nor2_1 _16832_ (.A(_08432_),
    .B(_10151_),
    .Y(_10237_));
 sky130_fd_sc_hd__a221o_1 _16833_ (.A1(\alu_shl[26] ),
    .A2(_10175_),
    .B1(_10123_),
    .B2(_08431_),
    .C1(_10237_),
    .X(_10238_));
 sky130_fd_sc_hd__a221o_1 _16834_ (.A1(\alu_shr[26] ),
    .A2(_10217_),
    .B1(_08434_),
    .B2(_10212_),
    .C1(_10227_),
    .X(_10239_));
 sky130_fd_sc_hd__o22a_1 _16835_ (.A1(net438),
    .A2(_10222_),
    .B1(_10238_),
    .B2(_10239_),
    .X(\alu_out[26] ));
 sky130_fd_sc_hd__clkbuf_2 _16836_ (.A(net286),
    .X(_10240_));
 sky130_fd_sc_hd__clkbuf_4 _16837_ (.A(_10240_),
    .X(_10241_));
 sky130_fd_sc_hd__a22o_1 _16838_ (.A1(\alu_shl[27] ),
    .A2(_10165_),
    .B1(_10113_),
    .B2(_08435_),
    .X(_10242_));
 sky130_fd_sc_hd__a31o_1 _16839_ (.A1(_10241_),
    .A2(_08436_),
    .A3(_10198_),
    .B1(_10242_),
    .X(_10243_));
 sky130_fd_sc_hd__a221o_1 _16840_ (.A1(\alu_shr[27] ),
    .A2(_10217_),
    .B1(_08439_),
    .B2(_10129_),
    .C1(_10227_),
    .X(_10244_));
 sky130_fd_sc_hd__o22a_1 _16841_ (.A1(net462),
    .A2(_10222_),
    .B1(_10243_),
    .B2(_10244_),
    .X(\alu_out[27] ));
 sky130_fd_sc_hd__clkbuf_2 _16842_ (.A(net287),
    .X(_10245_));
 sky130_fd_sc_hd__clkbuf_4 _16843_ (.A(_10245_),
    .X(_10246_));
 sky130_fd_sc_hd__a2bb2o_1 _16844_ (.A1_N(_08478_),
    .A2_N(_10150_),
    .B1(_10128_),
    .B2(\alu_shl[28] ),
    .X(_10247_));
 sky130_fd_sc_hd__a31o_1 _16845_ (.A1(_10246_),
    .A2(_08479_),
    .A3(_10198_),
    .B1(_10247_),
    .X(_10248_));
 sky130_fd_sc_hd__a221o_1 _16846_ (.A1(\alu_shr[28] ),
    .A2(_10095_),
    .B1(_08481_),
    .B2(_10129_),
    .C1(_10227_),
    .X(_10249_));
 sky130_fd_sc_hd__o22a_1 _16847_ (.A1(net422),
    .A2(_10222_),
    .B1(_10248_),
    .B2(_10249_),
    .X(\alu_out[28] ));
 sky130_fd_sc_hd__clkbuf_4 _16848_ (.A(_08397_),
    .X(_10250_));
 sky130_fd_sc_hd__a22o_1 _16849_ (.A1(\alu_shl[29] ),
    .A2(_10165_),
    .B1(_10113_),
    .B2(_08396_),
    .X(_10251_));
 sky130_fd_sc_hd__a31o_1 _16850_ (.A1(_10250_),
    .A2(_08398_),
    .A3(_10198_),
    .B1(_10251_),
    .X(_10252_));
 sky130_fd_sc_hd__a221o_1 _16851_ (.A1(\alu_shr[29] ),
    .A2(_10095_),
    .B1(_08400_),
    .B2(_10129_),
    .C1(_10227_),
    .X(_10253_));
 sky130_fd_sc_hd__o22a_1 _16852_ (.A1(net463),
    .A2(_10222_),
    .B1(_10252_),
    .B2(_10253_),
    .X(\alu_out[29] ));
 sky130_fd_sc_hd__clkbuf_2 _16853_ (.A(net290),
    .X(_10254_));
 sky130_fd_sc_hd__clkbuf_4 _16854_ (.A(_10254_),
    .X(_10255_));
 sky130_fd_sc_hd__a22o_1 _16855_ (.A1(\alu_shl[30] ),
    .A2(_10165_),
    .B1(_10113_),
    .B2(_08489_),
    .X(_10256_));
 sky130_fd_sc_hd__a31o_1 _16856_ (.A1(_10255_),
    .A2(_08487_),
    .A3(_10170_),
    .B1(_10256_),
    .X(_10257_));
 sky130_fd_sc_hd__a221o_1 _16857_ (.A1(\alu_shr[30] ),
    .A2(_10095_),
    .B1(_08490_),
    .B2(_10129_),
    .C1(_10093_),
    .X(_10258_));
 sky130_fd_sc_hd__o22a_1 _16858_ (.A1(\alu_add_sub[30] ),
    .A2(_10090_),
    .B1(_10257_),
    .B2(_10258_),
    .X(\alu_out[30] ));
 sky130_fd_sc_hd__clkbuf_4 _16859_ (.A(_08393_),
    .X(_10259_));
 sky130_fd_sc_hd__clkbuf_4 _16860_ (.A(net323),
    .X(_10260_));
 sky130_fd_sc_hd__a22o_1 _16861_ (.A1(\alu_shl[31] ),
    .A2(_10165_),
    .B1(_10113_),
    .B2(_08392_),
    .X(_10261_));
 sky130_fd_sc_hd__a31o_1 _16862_ (.A1(_10259_),
    .A2(_10260_),
    .A3(_10170_),
    .B1(_10261_),
    .X(_10262_));
 sky130_fd_sc_hd__a221o_1 _16863_ (.A1(\alu_shr[31] ),
    .A2(_10095_),
    .B1(_08395_),
    .B2(_10129_),
    .C1(_10093_),
    .X(_10263_));
 sky130_fd_sc_hd__o22a_1 _16864_ (.A1(net439),
    .A2(_10090_),
    .B1(_10262_),
    .B2(_10263_),
    .X(\alu_out[31] ));
 sky130_fd_sc_hd__clkbuf_4 _16865_ (.A(_08326_),
    .X(_10264_));
 sky130_fd_sc_hd__clkbuf_2 _16866_ (.A(_08677_),
    .X(_10265_));
 sky130_fd_sc_hd__a22o_2 _16867_ (.A1(_10264_),
    .A2(_08757_),
    .B1(_09213_),
    .B2(_10265_),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 _16868_ (.A(_09522_),
    .X(_10266_));
 sky130_vsdinv _16869_ (.A(_09213_),
    .Y(_10267_));
 sky130_fd_sc_hd__a211o_2 _16870_ (.A1(_08468_),
    .A2(_10104_),
    .B1(_10266_),
    .C1(_10267_),
    .X(net196));
 sky130_fd_sc_hd__a211o_2 _16871_ (.A1(_10264_),
    .A2(_10104_),
    .B1(_10266_),
    .C1(_10267_),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 _16872_ (.A(net161),
    .X(_10268_));
 sky130_fd_sc_hd__buf_2 _16873_ (.A(_10268_),
    .X(_10269_));
 sky130_fd_sc_hd__buf_4 _16874_ (.A(_10269_),
    .X(_10270_));
 sky130_fd_sc_hd__a22o_1 _16875_ (.A1(_10270_),
    .A2(_08511_),
    .B1(_10265_),
    .B2(_08484_),
    .X(net191));
 sky130_fd_sc_hd__a22o_1 _16876_ (.A1(_10108_),
    .A2(_08511_),
    .B1(_10265_),
    .B2(_10158_),
    .X(net192));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16877_ (.A(_08455_),
    .X(_10271_));
 sky130_fd_sc_hd__clkbuf_2 _16878_ (.A(_10271_),
    .X(_10272_));
 sky130_fd_sc_hd__buf_4 _16879_ (.A(_10272_),
    .X(_10273_));
 sky130_fd_sc_hd__a22o_2 _16880_ (.A1(_10273_),
    .A2(_08511_),
    .B1(_10265_),
    .B2(_10164_),
    .X(net162));
 sky130_fd_sc_hd__buf_2 _16881_ (.A(_08443_),
    .X(_10274_));
 sky130_fd_sc_hd__a22o_2 _16882_ (.A1(_10274_),
    .A2(_08511_),
    .B1(_10265_),
    .B2(_08413_),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_4 _16883_ (.A(net187),
    .X(_10275_));
 sky130_fd_sc_hd__clkbuf_2 _16884_ (.A(_10275_),
    .X(_10276_));
 sky130_fd_sc_hd__a22o_1 _16885_ (.A1(_10276_),
    .A2(_08511_),
    .B1(_10265_),
    .B2(_08343_),
    .X(net164));
 sky130_fd_sc_hd__buf_4 _16886_ (.A(net188),
    .X(_10277_));
 sky130_fd_sc_hd__clkbuf_2 _16887_ (.A(_08509_),
    .X(_10278_));
 sky130_fd_sc_hd__a22o_2 _16888_ (.A1(_10277_),
    .A2(_10278_),
    .B1(_08677_),
    .B2(_08347_),
    .X(net165));
 sky130_fd_sc_hd__buf_4 _16889_ (.A(net189),
    .X(_10279_));
 sky130_fd_sc_hd__a22o_2 _16890_ (.A1(_10279_),
    .A2(_10278_),
    .B1(_08677_),
    .B2(_08419_),
    .X(net166));
 sky130_fd_sc_hd__buf_4 _16891_ (.A(net190),
    .X(_10280_));
 sky130_fd_sc_hd__a22o_2 _16892_ (.A1(_10280_),
    .A2(_10278_),
    .B1(_08677_),
    .B2(_10188_),
    .X(net167));
 sky130_fd_sc_hd__buf_2 _16893_ (.A(_08469_),
    .X(_10281_));
 sky130_fd_sc_hd__buf_2 _16894_ (.A(_10281_),
    .X(_10282_));
 sky130_fd_sc_hd__mux2_1 _16895_ (.A0(_10282_),
    .A1(net306),
    .S(_09522_),
    .X(_10283_));
 sky130_fd_sc_hd__buf_1 _16896_ (.A(_10283_),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 _16897_ (.A(_10105_),
    .X(_10284_));
 sky130_fd_sc_hd__buf_2 _16898_ (.A(_10284_),
    .X(_10285_));
 sky130_fd_sc_hd__mux2_1 _16899_ (.A0(_10285_),
    .A1(_08383_),
    .S(_09522_),
    .X(_10286_));
 sky130_fd_sc_hd__buf_1 _16900_ (.A(_10286_),
    .X(net169));
 sky130_fd_sc_hd__buf_2 _16901_ (.A(_10271_),
    .X(_10287_));
 sky130_fd_sc_hd__clkbuf_4 _16902_ (.A(_08673_),
    .X(_10288_));
 sky130_fd_sc_hd__mux2_1 _16903_ (.A0(_10287_),
    .A1(net308),
    .S(_10288_),
    .X(_10289_));
 sky130_fd_sc_hd__buf_1 _16904_ (.A(_10289_),
    .X(net170));
 sky130_fd_sc_hd__mux2_1 _16905_ (.A0(_08443_),
    .A1(_08375_),
    .S(_10288_),
    .X(_10290_));
 sky130_fd_sc_hd__buf_1 _16906_ (.A(_10290_),
    .X(net171));
 sky130_fd_sc_hd__mux2_1 _16907_ (.A0(_10275_),
    .A1(net311),
    .S(_10288_),
    .X(_10291_));
 sky130_fd_sc_hd__clkbuf_2 _16908_ (.A(_10291_),
    .X(net173));
 sky130_fd_sc_hd__mux2_1 _16909_ (.A0(_10277_),
    .A1(_08364_),
    .S(_10288_),
    .X(_10292_));
 sky130_fd_sc_hd__buf_1 _16910_ (.A(_10292_),
    .X(net174));
 sky130_fd_sc_hd__mux2_1 _16911_ (.A0(_10279_),
    .A1(net313),
    .S(_10288_),
    .X(_10293_));
 sky130_fd_sc_hd__buf_1 _16912_ (.A(_10293_),
    .X(net175));
 sky130_fd_sc_hd__mux2_1 _16913_ (.A0(_10280_),
    .A1(_08369_),
    .S(_10288_),
    .X(_10294_));
 sky130_fd_sc_hd__clkbuf_2 _16914_ (.A(_10294_),
    .X(net176));
 sky130_fd_sc_hd__a22o_1 _16915_ (.A1(_08503_),
    .A2(_08484_),
    .B1(_10278_),
    .B2(_10270_),
    .X(_10295_));
 sky130_fd_sc_hd__a21o_1 _16916_ (.A1(net315),
    .A2(_10266_),
    .B1(_10295_),
    .X(net177));
 sky130_fd_sc_hd__a22o_1 _16917_ (.A1(_08503_),
    .A2(_10158_),
    .B1(_10278_),
    .B2(_10285_),
    .X(_10296_));
 sky130_fd_sc_hd__a21o_1 _16918_ (.A1(_08427_),
    .A2(_10266_),
    .B1(_10296_),
    .X(net178));
 sky130_fd_sc_hd__a22o_1 _16919_ (.A1(_08503_),
    .A2(_10164_),
    .B1(_10278_),
    .B2(_10287_),
    .X(_10297_));
 sky130_fd_sc_hd__a21o_1 _16920_ (.A1(net317),
    .A2(_10266_),
    .B1(_10297_),
    .X(net179));
 sky130_fd_sc_hd__buf_2 _16921_ (.A(_08443_),
    .X(_10298_));
 sky130_fd_sc_hd__a22o_1 _16922_ (.A1(_08503_),
    .A2(_08413_),
    .B1(_08510_),
    .B2(_10298_),
    .X(_10299_));
 sky130_fd_sc_hd__a21o_1 _16923_ (.A1(_08436_),
    .A2(_10266_),
    .B1(_10299_),
    .X(net180));
 sky130_fd_sc_hd__a22o_1 _16924_ (.A1(_08503_),
    .A2(_08343_),
    .B1(_08510_),
    .B2(_10275_),
    .X(_10300_));
 sky130_fd_sc_hd__a21o_2 _16925_ (.A1(_08479_),
    .A2(_09717_),
    .B1(_10300_),
    .X(net181));
 sky130_fd_sc_hd__a22o_1 _16926_ (.A1(_08324_),
    .A2(_08347_),
    .B1(_08510_),
    .B2(_10277_),
    .X(_10301_));
 sky130_fd_sc_hd__a21o_1 _16927_ (.A1(_08398_),
    .A2(_09717_),
    .B1(_10301_),
    .X(net182));
 sky130_fd_sc_hd__a22o_1 _16928_ (.A1(_08324_),
    .A2(_08419_),
    .B1(_08510_),
    .B2(_10279_),
    .X(_10302_));
 sky130_fd_sc_hd__a21o_2 _16929_ (.A1(_08487_),
    .A2(_09717_),
    .B1(_10302_),
    .X(net184));
 sky130_fd_sc_hd__a22o_1 _16930_ (.A1(_08324_),
    .A2(_10188_),
    .B1(_08510_),
    .B2(_10280_),
    .X(_10303_));
 sky130_fd_sc_hd__a21o_1 _16931_ (.A1(_10260_),
    .A2(_09717_),
    .B1(_10303_),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_2 _16932_ (.A(\irq_state[1] ),
    .X(_10304_));
 sky130_fd_sc_hd__buf_2 _16933_ (.A(_10304_),
    .X(_10305_));
 sky130_vsdinv _16934_ (.A(_10305_),
    .Y(_10306_));
 sky130_fd_sc_hd__or3_1 _16935_ (.A(\cpu_state[0] ),
    .B(_08148_),
    .C(_08539_),
    .X(_10307_));
 sky130_fd_sc_hd__or2_1 _16936_ (.A(\irq_pending[2] ),
    .B(net23),
    .X(_10308_));
 sky130_fd_sc_hd__o311a_1 _16937_ (.A1(_10306_),
    .A2(\irq_mask[2] ),
    .A3(_10307_),
    .B1(_10308_),
    .C1(_08321_),
    .X(_10309_));
 sky130_fd_sc_hd__or4_1 _16938_ (.A(_08202_),
    .B(_08188_),
    .C(_08199_),
    .D(_10309_),
    .X(_10310_));
 sky130_fd_sc_hd__clkbuf_1 _16939_ (.A(_10310_),
    .X(_00036_));
 sky130_fd_sc_hd__clkbuf_4 _16940_ (.A(_08456_),
    .X(_10311_));
 sky130_fd_sc_hd__nand2_1 _16941_ (.A(latched_branch),
    .B(latched_store),
    .Y(_10312_));
 sky130_fd_sc_hd__clkbuf_2 _16942_ (.A(_10312_),
    .X(_10313_));
 sky130_fd_sc_hd__clkbuf_2 _16943_ (.A(_10313_),
    .X(_10314_));
 sky130_fd_sc_hd__buf_2 _16944_ (.A(_10314_),
    .X(_10315_));
 sky130_fd_sc_hd__buf_2 _16945_ (.A(latched_branch),
    .X(_10316_));
 sky130_fd_sc_hd__buf_2 _16946_ (.A(latched_store),
    .X(_10317_));
 sky130_fd_sc_hd__a21o_1 _16947_ (.A1(_10316_),
    .A2(_10317_),
    .B1(\reg_next_pc[2] ),
    .X(_10318_));
 sky130_fd_sc_hd__o21a_1 _16948_ (.A1(\reg_out[2] ),
    .A2(_10315_),
    .B1(_10318_),
    .X(_10319_));
 sky130_fd_sc_hd__clkbuf_4 _16949_ (.A(_08523_),
    .X(_10320_));
 sky130_fd_sc_hd__mux2_1 _16950_ (.A0(_10311_),
    .A1(_10319_),
    .S(_10320_),
    .X(_10321_));
 sky130_fd_sc_hd__buf_2 _16951_ (.A(_10321_),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_4 _16952_ (.A(_08441_),
    .X(_10322_));
 sky130_fd_sc_hd__and2_1 _16953_ (.A(_10316_),
    .B(_10317_),
    .X(_10323_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16954_ (.A(_10323_),
    .X(_10324_));
 sky130_fd_sc_hd__clkbuf_2 _16955_ (.A(_10324_),
    .X(_10325_));
 sky130_fd_sc_hd__clkbuf_2 _16956_ (.A(_10325_),
    .X(_10326_));
 sky130_fd_sc_hd__clkbuf_2 _16957_ (.A(_10326_),
    .X(_10327_));
 sky130_fd_sc_hd__clkbuf_2 _16958_ (.A(_10327_),
    .X(_10328_));
 sky130_fd_sc_hd__mux2_1 _16959_ (.A0(\reg_next_pc[3] ),
    .A1(\reg_out[3] ),
    .S(_10328_),
    .X(_10329_));
 sky130_fd_sc_hd__mux2_1 _16960_ (.A0(_10322_),
    .A1(_10329_),
    .S(_10320_),
    .X(_10330_));
 sky130_fd_sc_hd__clkbuf_2 _16961_ (.A(_10330_),
    .X(net153));
 sky130_fd_sc_hd__buf_4 _16962_ (.A(_08475_),
    .X(_10331_));
 sky130_fd_sc_hd__mux2_1 _16963_ (.A0(\reg_next_pc[4] ),
    .A1(\reg_out[4] ),
    .S(_10328_),
    .X(_10332_));
 sky130_fd_sc_hd__mux2_1 _16964_ (.A0(_10331_),
    .A1(_10332_),
    .S(_10320_),
    .X(_10333_));
 sky130_fd_sc_hd__buf_2 _16965_ (.A(_10333_),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_4 _16966_ (.A(_08449_),
    .X(_10334_));
 sky130_fd_sc_hd__mux2_1 _16967_ (.A0(\reg_next_pc[5] ),
    .A1(\reg_out[5] ),
    .S(_10328_),
    .X(_10335_));
 sky130_fd_sc_hd__mux2_1 _16968_ (.A0(_10334_),
    .A1(_10335_),
    .S(_10320_),
    .X(_10336_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16969_ (.A(_10336_),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 _16970_ (.A(_08407_),
    .X(_10337_));
 sky130_fd_sc_hd__mux2_1 _16971_ (.A0(\reg_next_pc[6] ),
    .A1(\reg_out[6] ),
    .S(_10328_),
    .X(_10338_));
 sky130_fd_sc_hd__mux2_1 _16972_ (.A0(_10337_),
    .A1(_10338_),
    .S(_10320_),
    .X(_10339_));
 sky130_fd_sc_hd__clkbuf_2 _16973_ (.A(_10339_),
    .X(net156));
 sky130_fd_sc_hd__mux2_2 _16974_ (.A0(\reg_next_pc[7] ),
    .A1(\reg_out[7] ),
    .S(_10328_),
    .X(_10340_));
 sky130_fd_sc_hd__clkbuf_4 _16975_ (.A(_08523_),
    .X(_10341_));
 sky130_fd_sc_hd__buf_2 _16976_ (.A(_10341_),
    .X(_10342_));
 sky130_fd_sc_hd__mux2_1 _16977_ (.A0(_08461_),
    .A1(_10340_),
    .S(_10342_),
    .X(_10343_));
 sky130_fd_sc_hd__clkbuf_2 _16978_ (.A(_10343_),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 _16979_ (.A(_08482_),
    .X(_10344_));
 sky130_fd_sc_hd__mux2_1 _16980_ (.A0(\reg_next_pc[8] ),
    .A1(\reg_out[8] ),
    .S(_10328_),
    .X(_10345_));
 sky130_fd_sc_hd__mux2_1 _16981_ (.A0(_10344_),
    .A1(_10345_),
    .S(_10342_),
    .X(_10346_));
 sky130_fd_sc_hd__clkbuf_4 _16982_ (.A(_10346_),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 _16983_ (.A(_10327_),
    .X(_10347_));
 sky130_fd_sc_hd__mux2_1 _16984_ (.A0(\reg_next_pc[9] ),
    .A1(\reg_out[9] ),
    .S(_10347_),
    .X(_10348_));
 sky130_fd_sc_hd__mux2_1 _16985_ (.A0(_10157_),
    .A1(_10348_),
    .S(_10342_),
    .X(_10349_));
 sky130_fd_sc_hd__buf_2 _16986_ (.A(_10349_),
    .X(net159));
 sky130_fd_sc_hd__mux2_1 _16987_ (.A0(\reg_next_pc[10] ),
    .A1(\reg_out[10] ),
    .S(_10347_),
    .X(_10350_));
 sky130_fd_sc_hd__mux2_1 _16988_ (.A0(_10163_),
    .A1(_10350_),
    .S(_10342_),
    .X(_10351_));
 sky130_fd_sc_hd__clkbuf_2 _16989_ (.A(_10351_),
    .X(net130));
 sky130_fd_sc_hd__mux2_1 _16990_ (.A0(\reg_next_pc[11] ),
    .A1(\reg_out[11] ),
    .S(_10347_),
    .X(_10352_));
 sky130_fd_sc_hd__mux2_1 _16991_ (.A0(_08412_),
    .A1(_10352_),
    .S(_10342_),
    .X(_10353_));
 sky130_fd_sc_hd__clkbuf_4 _16992_ (.A(_10353_),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_4 _16993_ (.A(_08342_),
    .X(_10354_));
 sky130_fd_sc_hd__mux2_1 _16994_ (.A0(\reg_next_pc[12] ),
    .A1(\reg_out[12] ),
    .S(_10347_),
    .X(_10355_));
 sky130_fd_sc_hd__mux2_1 _16995_ (.A0(_10354_),
    .A1(_10355_),
    .S(_10342_),
    .X(_10356_));
 sky130_fd_sc_hd__clkbuf_2 _16996_ (.A(_10356_),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_4 _16997_ (.A(_08346_),
    .X(_10357_));
 sky130_fd_sc_hd__mux2_1 _16998_ (.A0(\reg_next_pc[13] ),
    .A1(\reg_out[13] ),
    .S(_10347_),
    .X(_10358_));
 sky130_fd_sc_hd__clkbuf_2 _16999_ (.A(_10341_),
    .X(_10359_));
 sky130_fd_sc_hd__mux2_1 _17000_ (.A0(_10357_),
    .A1(_10358_),
    .S(_10359_),
    .X(_10360_));
 sky130_fd_sc_hd__clkbuf_2 _17001_ (.A(_10360_),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_4 _17002_ (.A(_08417_),
    .X(_10361_));
 sky130_fd_sc_hd__mux2_1 _17003_ (.A0(\reg_next_pc[14] ),
    .A1(\reg_out[14] ),
    .S(_10347_),
    .X(_10362_));
 sky130_fd_sc_hd__mux2_1 _17004_ (.A0(_10361_),
    .A1(_10362_),
    .S(_10359_),
    .X(_10363_));
 sky130_fd_sc_hd__buf_2 _17005_ (.A(_10363_),
    .X(net134));
 sky130_fd_sc_hd__buf_2 _17006_ (.A(_10327_),
    .X(_10364_));
 sky130_fd_sc_hd__mux2_1 _17007_ (.A0(\reg_next_pc[15] ),
    .A1(\reg_out[15] ),
    .S(_10364_),
    .X(_10365_));
 sky130_fd_sc_hd__mux2_1 _17008_ (.A0(_10187_),
    .A1(_10365_),
    .S(_10359_),
    .X(_10366_));
 sky130_fd_sc_hd__buf_2 _17009_ (.A(_10366_),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_4 _17010_ (.A(_08378_),
    .X(_10367_));
 sky130_fd_sc_hd__mux2_1 _17011_ (.A0(\reg_next_pc[16] ),
    .A1(\reg_out[16] ),
    .S(_10364_),
    .X(_10368_));
 sky130_fd_sc_hd__mux2_1 _17012_ (.A0(_10367_),
    .A1(_10368_),
    .S(_10359_),
    .X(_10369_));
 sky130_fd_sc_hd__buf_2 _17013_ (.A(_10369_),
    .X(net136));
 sky130_fd_sc_hd__mux2_1 _17014_ (.A0(\reg_next_pc[17] ),
    .A1(\reg_out[17] ),
    .S(_10364_),
    .X(_10370_));
 sky130_fd_sc_hd__mux2_1 _17015_ (.A0(_10197_),
    .A1(_10370_),
    .S(_10359_),
    .X(_10371_));
 sky130_fd_sc_hd__clkbuf_4 _17016_ (.A(_10371_),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_4 _17017_ (.A(_08351_),
    .X(_10372_));
 sky130_fd_sc_hd__mux2_1 _17018_ (.A0(\reg_next_pc[18] ),
    .A1(\reg_out[18] ),
    .S(_10364_),
    .X(_10373_));
 sky130_fd_sc_hd__mux2_1 _17019_ (.A0(_10372_),
    .A1(_10373_),
    .S(_10359_),
    .X(_10374_));
 sky130_fd_sc_hd__buf_2 _17020_ (.A(_10374_),
    .X(net138));
 sky130_fd_sc_hd__mux2_1 _17021_ (.A0(\reg_next_pc[19] ),
    .A1(\reg_out[19] ),
    .S(_10364_),
    .X(_10375_));
 sky130_fd_sc_hd__clkbuf_2 _17022_ (.A(_10341_),
    .X(_10376_));
 sky130_fd_sc_hd__mux2_1 _17023_ (.A0(_10206_),
    .A1(_10375_),
    .S(_10376_),
    .X(_10377_));
 sky130_fd_sc_hd__buf_2 _17024_ (.A(_10377_),
    .X(net139));
 sky130_fd_sc_hd__buf_4 _17025_ (.A(_08355_),
    .X(_10378_));
 sky130_fd_sc_hd__mux2_1 _17026_ (.A0(\reg_next_pc[20] ),
    .A1(\reg_out[20] ),
    .S(_10364_),
    .X(_10379_));
 sky130_fd_sc_hd__mux2_1 _17027_ (.A0(_10378_),
    .A1(_10379_),
    .S(_10376_),
    .X(_10380_));
 sky130_fd_sc_hd__buf_2 _17028_ (.A(_10380_),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_2 _17029_ (.A(_10327_),
    .X(_10381_));
 sky130_fd_sc_hd__mux2_1 _17030_ (.A0(\reg_next_pc[21] ),
    .A1(\reg_out[21] ),
    .S(_10381_),
    .X(_10382_));
 sky130_fd_sc_hd__mux2_1 _17031_ (.A0(_10214_),
    .A1(_10382_),
    .S(_10376_),
    .X(_10383_));
 sky130_fd_sc_hd__buf_2 _17032_ (.A(_10383_),
    .X(net141));
 sky130_fd_sc_hd__buf_4 _17033_ (.A(_08359_),
    .X(_10384_));
 sky130_fd_sc_hd__mux2_1 _17034_ (.A0(\reg_next_pc[22] ),
    .A1(\reg_out[22] ),
    .S(_10381_),
    .X(_10385_));
 sky130_fd_sc_hd__mux2_1 _17035_ (.A0(_10384_),
    .A1(_10385_),
    .S(_10376_),
    .X(_10386_));
 sky130_fd_sc_hd__buf_2 _17036_ (.A(_10386_),
    .X(net142));
 sky130_fd_sc_hd__mux2_1 _17037_ (.A0(\reg_next_pc[23] ),
    .A1(\reg_out[23] ),
    .S(_10381_),
    .X(_10387_));
 sky130_fd_sc_hd__mux2_1 _17038_ (.A0(_10224_),
    .A1(_10387_),
    .S(_10376_),
    .X(_10388_));
 sky130_fd_sc_hd__buf_2 _17039_ (.A(_10388_),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_4 _17040_ (.A(_08423_),
    .X(_10389_));
 sky130_fd_sc_hd__mux2_1 _17041_ (.A0(\reg_next_pc[24] ),
    .A1(\reg_out[24] ),
    .S(_10381_),
    .X(_10390_));
 sky130_fd_sc_hd__mux2_1 _17042_ (.A0(_10389_),
    .A1(_10390_),
    .S(_10376_),
    .X(_10391_));
 sky130_fd_sc_hd__buf_2 _17043_ (.A(_10391_),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_4 _17044_ (.A(_10232_),
    .X(_10392_));
 sky130_fd_sc_hd__mux2_1 _17045_ (.A0(\reg_next_pc[25] ),
    .A1(\reg_out[25] ),
    .S(_10381_),
    .X(_10393_));
 sky130_fd_sc_hd__clkbuf_2 _17046_ (.A(_10341_),
    .X(_10394_));
 sky130_fd_sc_hd__mux2_1 _17047_ (.A0(_10392_),
    .A1(_10393_),
    .S(_10394_),
    .X(_10395_));
 sky130_fd_sc_hd__clkbuf_4 _17048_ (.A(_10395_),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 _17049_ (.A(net285),
    .X(_10396_));
 sky130_fd_sc_hd__clkbuf_4 _17050_ (.A(_10396_),
    .X(_10397_));
 sky130_fd_sc_hd__mux2_1 _17051_ (.A0(\reg_next_pc[26] ),
    .A1(\reg_out[26] ),
    .S(_10381_),
    .X(_10398_));
 sky130_fd_sc_hd__mux2_1 _17052_ (.A0(_10397_),
    .A1(_10398_),
    .S(_10394_),
    .X(_10399_));
 sky130_fd_sc_hd__buf_2 _17053_ (.A(_10399_),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 _17054_ (.A(_10327_),
    .X(_10400_));
 sky130_fd_sc_hd__mux2_1 _17055_ (.A0(\reg_next_pc[27] ),
    .A1(\reg_out[27] ),
    .S(_10400_),
    .X(_10401_));
 sky130_fd_sc_hd__mux2_1 _17056_ (.A0(_10241_),
    .A1(_10401_),
    .S(_10394_),
    .X(_10402_));
 sky130_fd_sc_hd__clkbuf_4 _17057_ (.A(_10402_),
    .X(net147));
 sky130_fd_sc_hd__mux2_1 _17058_ (.A0(\reg_next_pc[28] ),
    .A1(\reg_out[28] ),
    .S(_10400_),
    .X(_10403_));
 sky130_fd_sc_hd__mux2_1 _17059_ (.A0(_10246_),
    .A1(_10403_),
    .S(_10394_),
    .X(_10404_));
 sky130_fd_sc_hd__clkbuf_4 _17060_ (.A(_10404_),
    .X(net148));
 sky130_fd_sc_hd__mux2_1 _17061_ (.A0(\reg_next_pc[29] ),
    .A1(\reg_out[29] ),
    .S(_10400_),
    .X(_10405_));
 sky130_fd_sc_hd__mux2_1 _17062_ (.A0(_10250_),
    .A1(_10405_),
    .S(_10394_),
    .X(_10406_));
 sky130_fd_sc_hd__clkbuf_4 _17063_ (.A(_10406_),
    .X(net149));
 sky130_fd_sc_hd__mux2_1 _17064_ (.A0(\reg_next_pc[30] ),
    .A1(\reg_out[30] ),
    .S(_10400_),
    .X(_10407_));
 sky130_fd_sc_hd__mux2_1 _17065_ (.A0(_10255_),
    .A1(_10407_),
    .S(_10394_),
    .X(_10408_));
 sky130_fd_sc_hd__clkbuf_4 _17066_ (.A(_10408_),
    .X(net151));
 sky130_fd_sc_hd__mux2_1 _17067_ (.A0(\reg_next_pc[31] ),
    .A1(\reg_out[31] ),
    .S(_10400_),
    .X(_10409_));
 sky130_fd_sc_hd__mux2_1 _17068_ (.A0(_08393_),
    .A1(_10409_),
    .S(_10341_),
    .X(_10410_));
 sky130_fd_sc_hd__clkbuf_2 _17069_ (.A(_10410_),
    .X(net152));
 sky130_vsdinv _17070_ (.A(instr_sub),
    .Y(_10411_));
 sky130_fd_sc_hd__clkbuf_4 _17071_ (.A(_10411_),
    .X(_10412_));
 sky130_fd_sc_hd__nand2_1 _17072_ (.A(_10412_),
    .B(_10270_),
    .Y(_10413_));
 sky130_fd_sc_hd__nand2_1 _17073_ (.A(_10270_),
    .B(_08467_),
    .Y(_10414_));
 sky130_fd_sc_hd__a21o_1 _17074_ (.A1(_08468_),
    .A2(net161),
    .B1(_08467_),
    .X(_10415_));
 sky130_fd_sc_hd__o21a_1 _17075_ (.A1(_10264_),
    .A2(_10414_),
    .B1(_10415_),
    .X(_10416_));
 sky130_fd_sc_hd__xnor2_1 _17076_ (.A(_10413_),
    .B(_10416_),
    .Y(_00011_));
 sky130_fd_sc_hd__o21ai_1 _17077_ (.A1(_08672_),
    .A2(net172),
    .B1(_10415_),
    .Y(_10417_));
 sky130_fd_sc_hd__a22o_1 _17078_ (.A1(net267),
    .A2(net161),
    .B1(net172),
    .B2(net278),
    .X(_10418_));
 sky130_fd_sc_hd__nand2_1 _17079_ (.A(_08465_),
    .B(_10418_),
    .Y(_10419_));
 sky130_fd_sc_hd__mux2_1 _17080_ (.A0(_10417_),
    .A1(_10419_),
    .S(_10412_),
    .X(_10420_));
 sky130_fd_sc_hd__xnor2_1 _17081_ (.A(_08458_),
    .B(_10420_),
    .Y(_00022_));
 sky130_fd_sc_hd__nand2_1 _17082_ (.A(_08442_),
    .B(_08444_),
    .Y(_10421_));
 sky130_fd_sc_hd__nand2_1 _17083_ (.A(_08454_),
    .B(_08457_),
    .Y(_10422_));
 sky130_fd_sc_hd__and2b_1 _17084_ (.A_N(_08455_),
    .B(_08456_),
    .X(_10423_));
 sky130_fd_sc_hd__a21oi_1 _17085_ (.A1(_10422_),
    .A2(_10417_),
    .B1(_10423_),
    .Y(_10424_));
 sky130_fd_sc_hd__a31o_1 _17086_ (.A1(_08465_),
    .A2(_08454_),
    .A3(_10418_),
    .B1(_10124_),
    .X(_10425_));
 sky130_fd_sc_hd__clkbuf_4 _17087_ (.A(_10411_),
    .X(_10426_));
 sky130_fd_sc_hd__mux2_1 _17088_ (.A0(_10424_),
    .A1(_10425_),
    .S(_10426_),
    .X(_10427_));
 sky130_fd_sc_hd__xnor2_1 _17089_ (.A(_10421_),
    .B(_10427_),
    .Y(_00025_));
 sky130_fd_sc_hd__nand2_1 _17090_ (.A(_08474_),
    .B(_08476_),
    .Y(_10428_));
 sky130_fd_sc_hd__buf_2 _17091_ (.A(instr_sub),
    .X(_10429_));
 sky130_fd_sc_hd__clkbuf_4 _17092_ (.A(_10429_),
    .X(_10430_));
 sky130_vsdinv _17093_ (.A(_08443_),
    .Y(_10431_));
 sky130_fd_sc_hd__nand2_1 _17094_ (.A(_10431_),
    .B(_08441_),
    .Y(_10432_));
 sky130_fd_sc_hd__o21ai_1 _17095_ (.A1(_08445_),
    .A2(_10424_),
    .B1(_10432_),
    .Y(_10433_));
 sky130_fd_sc_hd__a311o_1 _17096_ (.A1(_08465_),
    .A2(_08454_),
    .A3(_10418_),
    .B1(_10124_),
    .C1(_10130_),
    .X(_10434_));
 sky130_fd_sc_hd__clkbuf_4 _17097_ (.A(instr_sub),
    .X(_10435_));
 sky130_fd_sc_hd__a21oi_1 _17098_ (.A1(_08442_),
    .A2(_10434_),
    .B1(_10435_),
    .Y(_10436_));
 sky130_fd_sc_hd__a21oi_1 _17099_ (.A1(_10430_),
    .A2(_10433_),
    .B1(_10436_),
    .Y(_10437_));
 sky130_fd_sc_hd__xnor2_1 _17100_ (.A(_10428_),
    .B(_10437_),
    .Y(_00026_));
 sky130_fd_sc_hd__and2b_1 _17101_ (.A_N(net187),
    .B(_08475_),
    .X(_10438_));
 sky130_fd_sc_hd__a21oi_1 _17102_ (.A1(_10428_),
    .A2(_10433_),
    .B1(_10438_),
    .Y(_10439_));
 sky130_fd_sc_hd__a31o_1 _17103_ (.A1(_08474_),
    .A2(_08442_),
    .A3(_10434_),
    .B1(_10134_),
    .X(_10440_));
 sky130_fd_sc_hd__mux2_1 _17104_ (.A0(_10439_),
    .A1(_10440_),
    .S(_10412_),
    .X(_10441_));
 sky130_fd_sc_hd__xor2_1 _17105_ (.A(_08453_),
    .B(_10441_),
    .X(_00027_));
 sky130_vsdinv _17106_ (.A(_08449_),
    .Y(_10442_));
 sky130_fd_sc_hd__a21o_1 _17107_ (.A1(net188),
    .A2(_10442_),
    .B1(_10439_),
    .X(_10443_));
 sky130_fd_sc_hd__o21ai_1 _17108_ (.A1(net188),
    .A2(_10442_),
    .B1(_10443_),
    .Y(_10444_));
 sky130_fd_sc_hd__a21oi_1 _17109_ (.A1(_08450_),
    .A2(_10440_),
    .B1(_08452_),
    .Y(_10445_));
 sky130_fd_sc_hd__mux2_1 _17110_ (.A0(_10444_),
    .A1(_10445_),
    .S(_10426_),
    .X(_10446_));
 sky130_fd_sc_hd__xnor2_1 _17111_ (.A(_08410_),
    .B(_10446_),
    .Y(_00028_));
 sky130_fd_sc_hd__nand2_1 _17112_ (.A(_08408_),
    .B(_08409_),
    .Y(_10447_));
 sky130_fd_sc_hd__and2b_1 _17113_ (.A_N(net189),
    .B(_08407_),
    .X(_10448_));
 sky130_fd_sc_hd__a21o_1 _17114_ (.A1(_10447_),
    .A2(_10444_),
    .B1(_10448_),
    .X(_10449_));
 sky130_fd_sc_hd__a211o_1 _17115_ (.A1(_08450_),
    .A2(_10440_),
    .B1(_08452_),
    .C1(_10141_),
    .X(_10450_));
 sky130_fd_sc_hd__nand2_1 _17116_ (.A(_08408_),
    .B(_10450_),
    .Y(_10451_));
 sky130_fd_sc_hd__mux2_1 _17117_ (.A0(_10449_),
    .A1(_10451_),
    .S(_10426_),
    .X(_10452_));
 sky130_fd_sc_hd__xnor2_1 _17118_ (.A(_08464_),
    .B(_10452_),
    .Y(_00029_));
 sky130_fd_sc_hd__a31oi_1 _17119_ (.A1(_08408_),
    .A2(_10145_),
    .A3(_10450_),
    .B1(_08463_),
    .Y(_10453_));
 sky130_vsdinv _17120_ (.A(net190),
    .Y(_10454_));
 sky130_fd_sc_hd__o21a_1 _17121_ (.A1(_10454_),
    .A2(_08460_),
    .B1(_10449_),
    .X(_10455_));
 sky130_fd_sc_hd__a21o_1 _17122_ (.A1(_10454_),
    .A2(_08460_),
    .B1(_10455_),
    .X(_10456_));
 sky130_fd_sc_hd__clkbuf_4 _17123_ (.A(instr_sub),
    .X(_10457_));
 sky130_fd_sc_hd__mux2_1 _17124_ (.A0(_10453_),
    .A1(_10456_),
    .S(_10457_),
    .X(_10458_));
 sky130_fd_sc_hd__xnor2_1 _17125_ (.A(_08486_),
    .B(_10458_),
    .Y(_00030_));
 sky130_vsdinv _17126_ (.A(_08486_),
    .Y(_10459_));
 sky130_fd_sc_hd__and2b_1 _17127_ (.A_N(_08484_),
    .B(_08482_),
    .X(_10460_));
 sky130_fd_sc_hd__a21o_1 _17128_ (.A1(_10459_),
    .A2(_10456_),
    .B1(_10460_),
    .X(_10461_));
 sky130_fd_sc_hd__o21ba_1 _17129_ (.A1(_10459_),
    .A2(_10453_),
    .B1_N(_08483_),
    .X(_10462_));
 sky130_fd_sc_hd__mux2_1 _17130_ (.A0(_10461_),
    .A1(_10462_),
    .S(_10426_),
    .X(_10463_));
 sky130_fd_sc_hd__xnor2_1 _17131_ (.A(_08391_),
    .B(_10463_),
    .Y(_00031_));
 sky130_fd_sc_hd__or2b_1 _17132_ (.A(_10156_),
    .B_N(net330),
    .X(_10464_));
 sky130_fd_sc_hd__and2b_1 _17133_ (.A_N(_10158_),
    .B(_10156_),
    .X(_10465_));
 sky130_fd_sc_hd__a21oi_1 _17134_ (.A1(_10461_),
    .A2(_10464_),
    .B1(_10465_),
    .Y(_10466_));
 sky130_fd_sc_hd__o21a_1 _17135_ (.A1(_08389_),
    .A2(_10462_),
    .B1(_08390_),
    .X(_10467_));
 sky130_fd_sc_hd__nor2_1 _17136_ (.A(_10435_),
    .B(_10467_),
    .Y(_10468_));
 sky130_fd_sc_hd__a21oi_1 _17137_ (.A1(_10430_),
    .A2(_10466_),
    .B1(_10468_),
    .Y(_10469_));
 sky130_fd_sc_hd__xnor2_1 _17138_ (.A(_08404_),
    .B(_10469_),
    .Y(_00001_));
 sky130_fd_sc_hd__or2b_1 _17139_ (.A(_10164_),
    .B_N(_08401_),
    .X(_10470_));
 sky130_fd_sc_hd__o21ai_1 _17140_ (.A1(_08404_),
    .A2(_10466_),
    .B1(_10470_),
    .Y(_10471_));
 sky130_fd_sc_hd__a21bo_1 _17141_ (.A1(_08402_),
    .A2(_10467_),
    .B1_N(_08403_),
    .X(_10472_));
 sky130_fd_sc_hd__mux2_1 _17142_ (.A0(_10471_),
    .A1(_10472_),
    .S(_10426_),
    .X(_10473_));
 sky130_fd_sc_hd__xnor2_1 _17143_ (.A(_08416_),
    .B(_10473_),
    .Y(_00002_));
 sky130_fd_sc_hd__nand2_1 _17144_ (.A(net269),
    .B(net301),
    .Y(_10474_));
 sky130_fd_sc_hd__a21oi_1 _17145_ (.A1(_10474_),
    .A2(_10472_),
    .B1(_08415_),
    .Y(_10475_));
 sky130_fd_sc_hd__and2b_1 _17146_ (.A_N(net301),
    .B(_08411_),
    .X(_10476_));
 sky130_fd_sc_hd__or2b_1 _17147_ (.A(_08411_),
    .B_N(_08413_),
    .X(_10477_));
 sky130_fd_sc_hd__o21a_1 _17148_ (.A1(_10471_),
    .A2(_10476_),
    .B1(_10477_),
    .X(_10478_));
 sky130_fd_sc_hd__nand2_1 _17149_ (.A(_10429_),
    .B(_10478_),
    .Y(_10479_));
 sky130_fd_sc_hd__o21ai_1 _17150_ (.A1(_10430_),
    .A2(_10475_),
    .B1(_10479_),
    .Y(_10480_));
 sky130_fd_sc_hd__xnor2_1 _17151_ (.A(_08345_),
    .B(_10480_),
    .Y(_00003_));
 sky130_fd_sc_hd__a2111o_1 _17152_ (.A1(_10474_),
    .A2(_10472_),
    .B1(_08415_),
    .C1(_08341_),
    .D1(_08344_),
    .X(_10481_));
 sky130_fd_sc_hd__mux2_1 _17153_ (.A0(_10354_),
    .A1(_10481_),
    .S(_10411_),
    .X(_10482_));
 sky130_vsdinv _17154_ (.A(_10482_),
    .Y(_10483_));
 sky130_fd_sc_hd__o22a_1 _17155_ (.A1(_08345_),
    .A2(_10479_),
    .B1(_10483_),
    .B2(_08341_),
    .X(_10484_));
 sky130_fd_sc_hd__xor2_1 _17156_ (.A(_08350_),
    .B(_10484_),
    .X(_00004_));
 sky130_vsdinv _17157_ (.A(_08347_),
    .Y(_10485_));
 sky130_fd_sc_hd__nor2_1 _17158_ (.A(_08345_),
    .B(_08350_),
    .Y(_10486_));
 sky130_fd_sc_hd__nor3b_1 _17159_ (.A(_08343_),
    .B(_08350_),
    .C_N(_08342_),
    .Y(_10487_));
 sky130_fd_sc_hd__a221o_1 _17160_ (.A1(_08346_),
    .A2(_10485_),
    .B1(_10486_),
    .B2(_10478_),
    .C1(_10487_),
    .X(_10488_));
 sky130_fd_sc_hd__nor2_1 _17161_ (.A(_08341_),
    .B(_08349_),
    .Y(_10489_));
 sky130_fd_sc_hd__a21o_1 _17162_ (.A1(_10481_),
    .A2(_10489_),
    .B1(_08348_),
    .X(_10490_));
 sky130_fd_sc_hd__mux2_1 _17163_ (.A0(_10488_),
    .A1(_10490_),
    .S(_10426_),
    .X(_10491_));
 sky130_fd_sc_hd__xnor2_1 _17164_ (.A(_08421_),
    .B(_10491_),
    .Y(_00005_));
 sky130_vsdinv _17165_ (.A(_08421_),
    .Y(_10492_));
 sky130_fd_sc_hd__and2b_1 _17166_ (.A_N(_08419_),
    .B(_08417_),
    .X(_10493_));
 sky130_fd_sc_hd__a21oi_1 _17167_ (.A1(_10492_),
    .A2(_10488_),
    .B1(_10493_),
    .Y(_10494_));
 sky130_fd_sc_hd__o21ba_1 _17168_ (.A1(_10492_),
    .A2(_10490_),
    .B1_N(_08418_),
    .X(_10495_));
 sky130_vsdinv _17169_ (.A(_10495_),
    .Y(_10496_));
 sky130_fd_sc_hd__mux2_1 _17170_ (.A0(_10494_),
    .A1(_10496_),
    .S(_10412_),
    .X(_10497_));
 sky130_fd_sc_hd__xor2_1 _17171_ (.A(_08448_),
    .B(_10497_),
    .X(_00006_));
 sky130_fd_sc_hd__or2b_1 _17172_ (.A(net305),
    .B_N(_10186_),
    .X(_10498_));
 sky130_fd_sc_hd__and2b_1 _17173_ (.A_N(_10186_),
    .B(_10188_),
    .X(_10499_));
 sky130_fd_sc_hd__a21o_1 _17174_ (.A1(_10494_),
    .A2(_10498_),
    .B1(_10499_),
    .X(_10500_));
 sky130_fd_sc_hd__o21ai_1 _17175_ (.A1(_08446_),
    .A2(_10495_),
    .B1(_08447_),
    .Y(_10501_));
 sky130_fd_sc_hd__mux2_1 _17176_ (.A0(_10500_),
    .A1(_10501_),
    .S(_10412_),
    .X(_10502_));
 sky130_fd_sc_hd__xor2_1 _17177_ (.A(_08381_),
    .B(_10502_),
    .X(_00007_));
 sky130_fd_sc_hd__a21oi_1 _17178_ (.A1(_08381_),
    .A2(_10501_),
    .B1(_08379_),
    .Y(_10503_));
 sky130_fd_sc_hd__or2b_1 _17179_ (.A(net306),
    .B_N(_08378_),
    .X(_10504_));
 sky130_fd_sc_hd__o211a_1 _17180_ (.A1(_08381_),
    .A2(_10500_),
    .B1(_10504_),
    .C1(_10429_),
    .X(_10505_));
 sky130_fd_sc_hd__o21ba_1 _17181_ (.A1(_10435_),
    .A2(_10503_),
    .B1_N(_10505_),
    .X(_10506_));
 sky130_fd_sc_hd__xnor2_1 _17182_ (.A(_08386_),
    .B(_10506_),
    .Y(_00008_));
 sky130_fd_sc_hd__nor2_1 _17183_ (.A(net275),
    .B(net307),
    .Y(_10507_));
 sky130_fd_sc_hd__o21a_1 _17184_ (.A1(_10507_),
    .A2(_10503_),
    .B1(_08385_),
    .X(_10508_));
 sky130_fd_sc_hd__or2b_1 _17185_ (.A(_08383_),
    .B_N(_08382_),
    .X(_10509_));
 sky130_fd_sc_hd__o221ai_2 _17186_ (.A1(_08387_),
    .A2(_10500_),
    .B1(_10504_),
    .B2(_08386_),
    .C1(_10509_),
    .Y(_10510_));
 sky130_fd_sc_hd__mux2_1 _17187_ (.A0(_10508_),
    .A1(_10510_),
    .S(_10457_),
    .X(_10511_));
 sky130_fd_sc_hd__xnor2_1 _17188_ (.A(_08354_),
    .B(_10511_),
    .Y(_00009_));
 sky130_fd_sc_hd__or2b_1 _17189_ (.A(_08354_),
    .B_N(_10510_),
    .X(_10512_));
 sky130_fd_sc_hd__or2b_1 _17190_ (.A(net308),
    .B_N(_08351_),
    .X(_10513_));
 sky130_fd_sc_hd__o21ba_1 _17191_ (.A1(_08353_),
    .A2(_10508_),
    .B1_N(_08352_),
    .X(_10514_));
 sky130_fd_sc_hd__nor2_1 _17192_ (.A(_10429_),
    .B(_10514_),
    .Y(_10515_));
 sky130_fd_sc_hd__a31o_1 _17193_ (.A1(_10430_),
    .A2(_10512_),
    .A3(_10513_),
    .B1(_10515_),
    .X(_10516_));
 sky130_fd_sc_hd__xor2_1 _17194_ (.A(_08377_),
    .B(_10516_),
    .X(_00010_));
 sky130_fd_sc_hd__or2b_1 _17195_ (.A(_08375_),
    .B_N(_08374_),
    .X(_10517_));
 sky130_fd_sc_hd__o21a_1 _17196_ (.A1(_08377_),
    .A2(_10513_),
    .B1(_10517_),
    .X(_10518_));
 sky130_fd_sc_hd__o21ai_1 _17197_ (.A1(_08377_),
    .A2(_10512_),
    .B1(_10518_),
    .Y(_10519_));
 sky130_fd_sc_hd__o21a_1 _17198_ (.A1(_08373_),
    .A2(_10514_),
    .B1(_08376_),
    .X(_10520_));
 sky130_fd_sc_hd__mux2_1 _17199_ (.A0(_10519_),
    .A1(_10520_),
    .S(_10411_),
    .X(_10521_));
 sky130_fd_sc_hd__xnor2_1 _17200_ (.A(_08358_),
    .B(_10521_),
    .Y(_00012_));
 sky130_fd_sc_hd__or2b_1 _17201_ (.A(_08358_),
    .B_N(_10519_),
    .X(_10522_));
 sky130_fd_sc_hd__or2b_1 _17202_ (.A(net311),
    .B_N(_08355_),
    .X(_10523_));
 sky130_fd_sc_hd__o21ba_1 _17203_ (.A1(_08357_),
    .A2(_10520_),
    .B1_N(_08356_),
    .X(_10524_));
 sky130_fd_sc_hd__nor2_1 _17204_ (.A(_10429_),
    .B(_10524_),
    .Y(_10525_));
 sky130_fd_sc_hd__a31o_1 _17205_ (.A1(_10435_),
    .A2(_10522_),
    .A3(_10523_),
    .B1(_10525_),
    .X(_10526_));
 sky130_fd_sc_hd__xor2_1 _17206_ (.A(_08367_),
    .B(_10526_),
    .X(_00013_));
 sky130_fd_sc_hd__or2b_1 _17207_ (.A(_08364_),
    .B_N(_08363_),
    .X(_10527_));
 sky130_fd_sc_hd__o21ai_1 _17208_ (.A1(_08367_),
    .A2(_10523_),
    .B1(_10527_),
    .Y(_10528_));
 sky130_fd_sc_hd__o21bai_1 _17209_ (.A1(_08367_),
    .A2(_10522_),
    .B1_N(_10528_),
    .Y(_10529_));
 sky130_fd_sc_hd__o21a_1 _17210_ (.A1(_08365_),
    .A2(_10524_),
    .B1(_08366_),
    .X(_10530_));
 sky130_fd_sc_hd__mux2_1 _17211_ (.A0(_10529_),
    .A1(_10530_),
    .S(_10411_),
    .X(_10531_));
 sky130_fd_sc_hd__xnor2_1 _17212_ (.A(_08362_),
    .B(_10531_),
    .Y(_00014_));
 sky130_fd_sc_hd__or2_1 _17213_ (.A(_08360_),
    .B(_08361_),
    .X(_10532_));
 sky130_fd_sc_hd__o21ba_1 _17214_ (.A1(_10532_),
    .A2(_10530_),
    .B1_N(_08360_),
    .X(_10533_));
 sky130_fd_sc_hd__and2b_1 _17215_ (.A_N(net313),
    .B(_08359_),
    .X(_10534_));
 sky130_fd_sc_hd__a21o_1 _17216_ (.A1(_10532_),
    .A2(_10529_),
    .B1(_10534_),
    .X(_10535_));
 sky130_fd_sc_hd__mux2_1 _17217_ (.A0(_10533_),
    .A1(_10535_),
    .S(_10457_),
    .X(_10536_));
 sky130_fd_sc_hd__xnor2_1 _17218_ (.A(_08371_),
    .B(_10536_),
    .Y(_00015_));
 sky130_fd_sc_hd__a21oi_1 _17219_ (.A1(_10532_),
    .A2(_10528_),
    .B1(_10534_),
    .Y(_10537_));
 sky130_fd_sc_hd__or2b_1 _17220_ (.A(_08369_),
    .B_N(_10223_),
    .X(_10538_));
 sky130_fd_sc_hd__o221a_1 _17221_ (.A1(_08372_),
    .A2(_10518_),
    .B1(_10537_),
    .B2(_08371_),
    .C1(_10538_),
    .X(_10539_));
 sky130_fd_sc_hd__o31a_1 _17222_ (.A1(_08372_),
    .A2(_08377_),
    .A3(_10512_),
    .B1(_10539_),
    .X(_10540_));
 sky130_fd_sc_hd__a21oi_1 _17223_ (.A1(_08370_),
    .A2(_10533_),
    .B1(_08368_),
    .Y(_10541_));
 sky130_fd_sc_hd__mux2_1 _17224_ (.A0(_10540_),
    .A1(_10541_),
    .S(_10412_),
    .X(_10542_));
 sky130_fd_sc_hd__xor2_1 _17225_ (.A(_08426_),
    .B(_10542_),
    .X(_00016_));
 sky130_fd_sc_hd__a21o_1 _17226_ (.A1(_08426_),
    .A2(_10541_),
    .B1(_08424_),
    .X(_10543_));
 sky130_fd_sc_hd__or2b_1 _17227_ (.A(net315),
    .B_N(_08423_),
    .X(_10544_));
 sky130_fd_sc_hd__o21a_1 _17228_ (.A1(_08426_),
    .A2(_10540_),
    .B1(_10544_),
    .X(_10545_));
 sky130_fd_sc_hd__mux2_1 _17229_ (.A0(_10543_),
    .A1(_10545_),
    .S(_10435_),
    .X(_10546_));
 sky130_fd_sc_hd__xor2_1 _17230_ (.A(_08430_),
    .B(_10546_),
    .X(_00017_));
 sky130_fd_sc_hd__a21oi_1 _17231_ (.A1(_10233_),
    .A2(_10543_),
    .B1(_08429_),
    .Y(_10547_));
 sky130_fd_sc_hd__or2b_1 _17232_ (.A(_08427_),
    .B_N(_10232_),
    .X(_10548_));
 sky130_fd_sc_hd__o21ai_1 _17233_ (.A1(_08430_),
    .A2(_10544_),
    .B1(_10548_),
    .Y(_10549_));
 sky130_fd_sc_hd__nor3_1 _17234_ (.A(_08426_),
    .B(_08430_),
    .C(_10540_),
    .Y(_10550_));
 sky130_fd_sc_hd__or2_1 _17235_ (.A(_10549_),
    .B(_10550_),
    .X(_10551_));
 sky130_fd_sc_hd__mux2_1 _17236_ (.A0(_10547_),
    .A1(_10551_),
    .S(_10457_),
    .X(_10552_));
 sky130_fd_sc_hd__xnor2_1 _17237_ (.A(_08434_),
    .B(_10552_),
    .Y(_00018_));
 sky130_fd_sc_hd__o21bai_1 _17238_ (.A1(_08433_),
    .A2(_10547_),
    .B1_N(_08431_),
    .Y(_10553_));
 sky130_fd_sc_hd__and2b_1 _17239_ (.A_N(net317),
    .B(_10396_),
    .X(_10554_));
 sky130_fd_sc_hd__a21oi_1 _17240_ (.A1(_08433_),
    .A2(_10551_),
    .B1(_10554_),
    .Y(_10555_));
 sky130_fd_sc_hd__mux2_1 _17241_ (.A0(_10553_),
    .A1(_10555_),
    .S(_10457_),
    .X(_10556_));
 sky130_fd_sc_hd__xnor2_1 _17242_ (.A(_08438_),
    .B(_10556_),
    .Y(_00019_));
 sky130_fd_sc_hd__a21boi_1 _17243_ (.A1(_08435_),
    .A2(_10553_),
    .B1_N(_08437_),
    .Y(_10557_));
 sky130_fd_sc_hd__a21o_1 _17244_ (.A1(_08433_),
    .A2(_10549_),
    .B1(_10554_),
    .X(_10558_));
 sky130_vsdinv _17245_ (.A(_08436_),
    .Y(_10559_));
 sky130_fd_sc_hd__a2bb2o_1 _17246_ (.A1_N(_10540_),
    .A2_N(_08440_),
    .B1(_10559_),
    .B2(_10240_),
    .X(_10560_));
 sky130_fd_sc_hd__a21o_1 _17247_ (.A1(_08438_),
    .A2(_10558_),
    .B1(_10560_),
    .X(_10561_));
 sky130_fd_sc_hd__mux2_1 _17248_ (.A0(_10557_),
    .A1(_10561_),
    .S(_10457_),
    .X(_10562_));
 sky130_fd_sc_hd__xnor2_1 _17249_ (.A(_08481_),
    .B(_10562_),
    .Y(_00020_));
 sky130_fd_sc_hd__o21ai_1 _17250_ (.A1(_08478_),
    .A2(_10557_),
    .B1(_08480_),
    .Y(_10563_));
 sky130_vsdinv _17251_ (.A(_08481_),
    .Y(_10564_));
 sky130_fd_sc_hd__and2b_1 _17252_ (.A_N(_08479_),
    .B(_10245_),
    .X(_10565_));
 sky130_fd_sc_hd__a21oi_1 _17253_ (.A1(_10564_),
    .A2(_10561_),
    .B1(_10565_),
    .Y(_10566_));
 sky130_fd_sc_hd__mux2_1 _17254_ (.A0(_10563_),
    .A1(_10566_),
    .S(_10435_),
    .X(_10567_));
 sky130_fd_sc_hd__xor2_1 _17255_ (.A(_08400_),
    .B(_10567_),
    .X(_00021_));
 sky130_fd_sc_hd__nand2_1 _17256_ (.A(_08488_),
    .B(_08489_),
    .Y(_10568_));
 sky130_fd_sc_hd__or2b_1 _17257_ (.A(net320),
    .B_N(_08397_),
    .X(_10569_));
 sky130_fd_sc_hd__and2b_1 _17258_ (.A_N(_08397_),
    .B(_08398_),
    .X(_10570_));
 sky130_fd_sc_hd__a21oi_1 _17259_ (.A1(_10566_),
    .A2(_10569_),
    .B1(_10570_),
    .Y(_10571_));
 sky130_fd_sc_hd__a21oi_1 _17260_ (.A1(_08396_),
    .A2(_10563_),
    .B1(instr_sub),
    .Y(_10572_));
 sky130_fd_sc_hd__and2_1 _17261_ (.A(_08399_),
    .B(_10572_),
    .X(_10573_));
 sky130_fd_sc_hd__a21oi_1 _17262_ (.A1(_10430_),
    .A2(_10571_),
    .B1(_10573_),
    .Y(_10574_));
 sky130_fd_sc_hd__xnor2_1 _17263_ (.A(_10568_),
    .B(_10574_),
    .Y(_00023_));
 sky130_fd_sc_hd__a21bo_1 _17264_ (.A1(_10429_),
    .A2(_10255_),
    .B1_N(_08489_),
    .X(_10575_));
 sky130_fd_sc_hd__or2b_1 _17265_ (.A(_08487_),
    .B_N(_10255_),
    .X(_10576_));
 sky130_fd_sc_hd__or3b_1 _17266_ (.A(_10411_),
    .B(_10571_),
    .C_N(_10576_),
    .X(_10577_));
 sky130_fd_sc_hd__a22o_1 _17267_ (.A1(_08488_),
    .A2(_10573_),
    .B1(_10575_),
    .B2(_10577_),
    .X(_10578_));
 sky130_fd_sc_hd__xnor2_1 _17268_ (.A(_08395_),
    .B(_10578_),
    .Y(_00024_));
 sky130_fd_sc_hd__or2b_1 _17269_ (.A(net323),
    .B_N(_10259_),
    .X(_10579_));
 sky130_fd_sc_hd__nand2_1 _17270_ (.A(_10568_),
    .B(_10571_),
    .Y(_10580_));
 sky130_fd_sc_hd__and2b_1 _17271_ (.A_N(_10259_),
    .B(_10260_),
    .X(_10581_));
 sky130_fd_sc_hd__a31o_1 _17272_ (.A1(_10576_),
    .A2(_10579_),
    .A3(_10580_),
    .B1(_10581_),
    .X(_00034_));
 sky130_fd_sc_hd__o21ba_1 _17273_ (.A1(_08395_),
    .A2(_00034_),
    .B1_N(_10581_),
    .X(_00033_));
 sky130_fd_sc_hd__buf_2 _17274_ (.A(\genblk1.pcpi_mul.rs2[0] ),
    .X(_10582_));
 sky130_fd_sc_hd__clkbuf_2 _17275_ (.A(_10582_),
    .X(_10583_));
 sky130_fd_sc_hd__clkbuf_4 _17276_ (.A(_10583_),
    .X(_10584_));
 sky130_fd_sc_hd__buf_2 _17277_ (.A(_10584_),
    .X(_10585_));
 sky130_fd_sc_hd__clkbuf_4 _17278_ (.A(_10585_),
    .X(_10586_));
 sky130_fd_sc_hd__clkbuf_2 _17279_ (.A(\genblk1.pcpi_mul.rs1[0] ),
    .X(_10587_));
 sky130_fd_sc_hd__clkbuf_2 _17280_ (.A(_10587_),
    .X(_10588_));
 sky130_fd_sc_hd__buf_2 _17281_ (.A(_10588_),
    .X(_10589_));
 sky130_fd_sc_hd__clkbuf_4 _17282_ (.A(_10589_),
    .X(_10590_));
 sky130_fd_sc_hd__buf_2 _17283_ (.A(_10590_),
    .X(_10591_));
 sky130_fd_sc_hd__buf_2 _17284_ (.A(_10591_),
    .X(_10592_));
 sky130_fd_sc_hd__and2_1 _17285_ (.A(_10586_),
    .B(_10592_),
    .X(_10593_));
 sky130_fd_sc_hd__clkbuf_1 _17286_ (.A(_10593_),
    .X(_00050_));
 sky130_fd_sc_hd__buf_2 _17287_ (.A(\genblk1.pcpi_mul.rs1[1] ),
    .X(_10594_));
 sky130_fd_sc_hd__clkbuf_2 _17288_ (.A(_10594_),
    .X(_10595_));
 sky130_fd_sc_hd__clkbuf_4 _17289_ (.A(_10595_),
    .X(_10596_));
 sky130_fd_sc_hd__buf_2 _17290_ (.A(_10596_),
    .X(_10597_));
 sky130_fd_sc_hd__clkbuf_4 _17291_ (.A(_10597_),
    .X(_10598_));
 sky130_fd_sc_hd__buf_2 _17292_ (.A(\genblk1.pcpi_mul.rs2[1] ),
    .X(_10599_));
 sky130_fd_sc_hd__buf_4 _17293_ (.A(_10599_),
    .X(_10600_));
 sky130_fd_sc_hd__buf_2 _17294_ (.A(_10600_),
    .X(_10601_));
 sky130_fd_sc_hd__clkbuf_2 _17295_ (.A(_10601_),
    .X(_10602_));
 sky130_fd_sc_hd__buf_2 _17296_ (.A(_10592_),
    .X(_10603_));
 sky130_fd_sc_hd__a22oi_1 _17297_ (.A1(_10586_),
    .A2(_10598_),
    .B1(_10602_),
    .B2(_10603_),
    .Y(_10604_));
 sky130_fd_sc_hd__and3_1 _17298_ (.A(_10598_),
    .B(_10602_),
    .C(_00050_),
    .X(_10605_));
 sky130_fd_sc_hd__nor2_1 _17299_ (.A(_10604_),
    .B(_10605_),
    .Y(_00051_));
 sky130_fd_sc_hd__clkbuf_2 _17300_ (.A(\genblk1.pcpi_mul.rs1[2] ),
    .X(_10606_));
 sky130_fd_sc_hd__buf_2 _17301_ (.A(_10606_),
    .X(_10607_));
 sky130_fd_sc_hd__clkbuf_4 _17302_ (.A(_10607_),
    .X(_10608_));
 sky130_fd_sc_hd__buf_4 _17303_ (.A(_10608_),
    .X(_10609_));
 sky130_fd_sc_hd__buf_2 _17304_ (.A(\genblk1.pcpi_mul.rs2[2] ),
    .X(_10610_));
 sky130_fd_sc_hd__buf_4 _17305_ (.A(_10610_),
    .X(_10611_));
 sky130_fd_sc_hd__buf_2 _17306_ (.A(_10611_),
    .X(_10612_));
 sky130_fd_sc_hd__buf_4 _17307_ (.A(_10612_),
    .X(_10613_));
 sky130_fd_sc_hd__a22o_1 _17308_ (.A1(_10597_),
    .A2(_10602_),
    .B1(_10613_),
    .B2(_10591_),
    .X(_10614_));
 sky130_fd_sc_hd__and4_1 _17309_ (.A(_10590_),
    .B(_10597_),
    .C(_10602_),
    .D(_10613_),
    .X(_10615_));
 sky130_vsdinv _17310_ (.A(_10615_),
    .Y(_10616_));
 sky130_fd_sc_hd__and4_1 _17311_ (.A(_10586_),
    .B(_10609_),
    .C(_10614_),
    .D(_10616_),
    .X(_10617_));
 sky130_fd_sc_hd__a22oi_1 _17312_ (.A1(_10586_),
    .A2(_10609_),
    .B1(_10614_),
    .B2(_10616_),
    .Y(_10618_));
 sky130_fd_sc_hd__nor2_1 _17313_ (.A(_10617_),
    .B(_10618_),
    .Y(_10619_));
 sky130_fd_sc_hd__nand2_1 _17314_ (.A(_10605_),
    .B(_10619_),
    .Y(_10620_));
 sky130_fd_sc_hd__or2_1 _17315_ (.A(_10605_),
    .B(_10619_),
    .X(_10621_));
 sky130_fd_sc_hd__and2_1 _17316_ (.A(_10620_),
    .B(_10621_),
    .X(_10622_));
 sky130_fd_sc_hd__clkbuf_1 _17317_ (.A(_10622_),
    .X(_00052_));
 sky130_fd_sc_hd__buf_2 _17318_ (.A(_10589_),
    .X(_10623_));
 sky130_fd_sc_hd__buf_2 _17319_ (.A(\genblk1.pcpi_mul.rs2[3] ),
    .X(_10624_));
 sky130_fd_sc_hd__clkbuf_4 _17320_ (.A(_10624_),
    .X(_10625_));
 sky130_fd_sc_hd__buf_2 _17321_ (.A(_10625_),
    .X(_10626_));
 sky130_fd_sc_hd__clkbuf_2 _17322_ (.A(_10600_),
    .X(_10627_));
 sky130_fd_sc_hd__buf_2 _17323_ (.A(\genblk1.pcpi_mul.rs1[2] ),
    .X(_10628_));
 sky130_fd_sc_hd__buf_1 _17324_ (.A(_10628_),
    .X(_10629_));
 sky130_fd_sc_hd__buf_2 _17325_ (.A(_10629_),
    .X(_10630_));
 sky130_fd_sc_hd__buf_2 _17326_ (.A(\genblk1.pcpi_mul.rs2[2] ),
    .X(_10631_));
 sky130_fd_sc_hd__clkbuf_2 _17327_ (.A(_10631_),
    .X(_10632_));
 sky130_fd_sc_hd__clkbuf_2 _17328_ (.A(_10632_),
    .X(_10633_));
 sky130_fd_sc_hd__clkbuf_2 _17329_ (.A(\genblk1.pcpi_mul.rs1[1] ),
    .X(_10634_));
 sky130_fd_sc_hd__clkbuf_2 _17330_ (.A(_10634_),
    .X(_10635_));
 sky130_fd_sc_hd__clkbuf_4 _17331_ (.A(_10635_),
    .X(_10636_));
 sky130_fd_sc_hd__a22oi_1 _17332_ (.A1(_10627_),
    .A2(_10630_),
    .B1(_10633_),
    .B2(_10636_),
    .Y(_10637_));
 sky130_fd_sc_hd__clkbuf_2 _17333_ (.A(_10635_),
    .X(_10638_));
 sky130_fd_sc_hd__buf_2 _17334_ (.A(\genblk1.pcpi_mul.rs2[1] ),
    .X(_10639_));
 sky130_fd_sc_hd__clkbuf_4 _17335_ (.A(_10639_),
    .X(_10640_));
 sky130_fd_sc_hd__buf_2 _17336_ (.A(_10640_),
    .X(_10641_));
 sky130_fd_sc_hd__and4_1 _17337_ (.A(_10638_),
    .B(_10641_),
    .C(_10608_),
    .D(_10632_),
    .X(_10642_));
 sky130_fd_sc_hd__o2bb2a_1 _17338_ (.A1_N(_10623_),
    .A2_N(_10626_),
    .B1(_10637_),
    .B2(_10642_),
    .X(_10643_));
 sky130_fd_sc_hd__clkbuf_4 _17339_ (.A(\genblk1.pcpi_mul.rs2[3] ),
    .X(_10644_));
 sky130_fd_sc_hd__clkbuf_2 _17340_ (.A(_10644_),
    .X(_10645_));
 sky130_fd_sc_hd__and4bb_1 _17341_ (.A_N(_10637_),
    .B_N(_10642_),
    .C(_10623_),
    .D(_10645_),
    .X(_10646_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17342_ (.A(\genblk1.pcpi_mul.rs1[3] ),
    .X(_10647_));
 sky130_fd_sc_hd__clkbuf_2 _17343_ (.A(_10647_),
    .X(_10648_));
 sky130_fd_sc_hd__buf_2 _17344_ (.A(_10648_),
    .X(_10649_));
 sky130_fd_sc_hd__buf_2 _17345_ (.A(_10649_),
    .X(_10650_));
 sky130_fd_sc_hd__clkbuf_4 _17346_ (.A(_10650_),
    .X(_10651_));
 sky130_fd_sc_hd__and4bb_1 _17347_ (.A_N(_10643_),
    .B_N(_10646_),
    .C(_10585_),
    .D(_10651_),
    .X(_10652_));
 sky130_fd_sc_hd__o2bb2a_1 _17348_ (.A1_N(_10585_),
    .A2_N(_10651_),
    .B1(_10643_),
    .B2(_10646_),
    .X(_10653_));
 sky130_fd_sc_hd__nor2_1 _17349_ (.A(_10652_),
    .B(_10653_),
    .Y(_10654_));
 sky130_fd_sc_hd__nand2_1 _17350_ (.A(_10617_),
    .B(_10654_),
    .Y(_10655_));
 sky130_fd_sc_hd__or2_1 _17351_ (.A(_10617_),
    .B(_10654_),
    .X(_10656_));
 sky130_fd_sc_hd__a21oi_1 _17352_ (.A1(_10655_),
    .A2(_10656_),
    .B1(_10615_),
    .Y(_10657_));
 sky130_fd_sc_hd__a21o_1 _17353_ (.A1(_10615_),
    .A2(_10654_),
    .B1(_10657_),
    .X(_10658_));
 sky130_fd_sc_hd__nor2_1 _17354_ (.A(_10620_),
    .B(_10658_),
    .Y(_10659_));
 sky130_fd_sc_hd__and2_1 _17355_ (.A(_10620_),
    .B(_10658_),
    .X(_10660_));
 sky130_fd_sc_hd__nor2_1 _17356_ (.A(_10659_),
    .B(_10660_),
    .Y(_00053_));
 sky130_fd_sc_hd__clkbuf_2 _17357_ (.A(\genblk1.pcpi_mul.rs2[4] ),
    .X(_10661_));
 sky130_fd_sc_hd__buf_2 _17358_ (.A(_10661_),
    .X(_10662_));
 sky130_fd_sc_hd__clkbuf_8 _17359_ (.A(_10662_),
    .X(_10663_));
 sky130_fd_sc_hd__clkbuf_2 _17360_ (.A(\genblk1.pcpi_mul.rs1[4] ),
    .X(_10664_));
 sky130_fd_sc_hd__clkbuf_2 _17361_ (.A(_10664_),
    .X(_10665_));
 sky130_fd_sc_hd__buf_2 _17362_ (.A(_10665_),
    .X(_10666_));
 sky130_fd_sc_hd__clkbuf_4 _17363_ (.A(_10666_),
    .X(_10667_));
 sky130_fd_sc_hd__a22oi_1 _17364_ (.A1(_10623_),
    .A2(_10663_),
    .B1(_10667_),
    .B2(_10584_),
    .Y(_10668_));
 sky130_fd_sc_hd__buf_2 _17365_ (.A(_10582_),
    .X(_10669_));
 sky130_fd_sc_hd__clkbuf_2 _17366_ (.A(\genblk1.pcpi_mul.rs2[4] ),
    .X(_10670_));
 sky130_fd_sc_hd__clkbuf_4 _17367_ (.A(_10670_),
    .X(_10671_));
 sky130_fd_sc_hd__buf_2 _17368_ (.A(_10671_),
    .X(_10672_));
 sky130_fd_sc_hd__and4_2 _17369_ (.A(_10669_),
    .B(_10588_),
    .C(_10672_),
    .D(_10666_),
    .X(_10673_));
 sky130_fd_sc_hd__nor2_1 _17370_ (.A(_10668_),
    .B(_10673_),
    .Y(_10674_));
 sky130_fd_sc_hd__buf_2 _17371_ (.A(_10648_),
    .X(_10675_));
 sky130_fd_sc_hd__clkbuf_4 _17372_ (.A(_10675_),
    .X(_10676_));
 sky130_fd_sc_hd__a22o_1 _17373_ (.A1(_10630_),
    .A2(_10633_),
    .B1(_10676_),
    .B2(_10601_),
    .X(_10677_));
 sky130_fd_sc_hd__nand4_1 _17374_ (.A(_10601_),
    .B(_10630_),
    .C(_10633_),
    .D(_10651_),
    .Y(_10678_));
 sky130_fd_sc_hd__a22o_1 _17375_ (.A1(_10596_),
    .A2(_10626_),
    .B1(_10677_),
    .B2(_10678_),
    .X(_10679_));
 sky130_fd_sc_hd__buf_2 _17376_ (.A(_10645_),
    .X(_10680_));
 sky130_fd_sc_hd__nand4_1 _17377_ (.A(_10597_),
    .B(_10680_),
    .C(_10677_),
    .D(_10678_),
    .Y(_10681_));
 sky130_fd_sc_hd__nand3_1 _17378_ (.A(_10674_),
    .B(_10679_),
    .C(_10681_),
    .Y(_10682_));
 sky130_fd_sc_hd__a21o_1 _17379_ (.A1(_10679_),
    .A2(_10681_),
    .B1(_10674_),
    .X(_10683_));
 sky130_fd_sc_hd__and3_1 _17380_ (.A(_10652_),
    .B(_10682_),
    .C(_10683_),
    .X(_10684_));
 sky130_fd_sc_hd__a21oi_1 _17381_ (.A1(_10682_),
    .A2(_10683_),
    .B1(_10652_),
    .Y(_10685_));
 sky130_fd_sc_hd__nor2_1 _17382_ (.A(_10684_),
    .B(_10685_),
    .Y(_10686_));
 sky130_fd_sc_hd__nor2_1 _17383_ (.A(_10642_),
    .B(_10646_),
    .Y(_10687_));
 sky130_fd_sc_hd__xnor2_1 _17384_ (.A(_10686_),
    .B(_10687_),
    .Y(_10688_));
 sky130_fd_sc_hd__o21a_1 _17385_ (.A1(_10615_),
    .A2(_10617_),
    .B1(_10654_),
    .X(_10689_));
 sky130_fd_sc_hd__and2_1 _17386_ (.A(_10688_),
    .B(_10689_),
    .X(_10690_));
 sky130_fd_sc_hd__or2_1 _17387_ (.A(_10688_),
    .B(_10689_),
    .X(_10691_));
 sky130_fd_sc_hd__or2b_1 _17388_ (.A(_10690_),
    .B_N(_10691_),
    .X(_10692_));
 sky130_fd_sc_hd__xnor2_1 _17389_ (.A(_10659_),
    .B(_10692_),
    .Y(_00054_));
 sky130_fd_sc_hd__o21bai_1 _17390_ (.A1(_10685_),
    .A2(_10687_),
    .B1_N(_10684_),
    .Y(_10693_));
 sky130_fd_sc_hd__nand2_1 _17391_ (.A(_10678_),
    .B(_10681_),
    .Y(_10694_));
 sky130_fd_sc_hd__clkbuf_4 _17392_ (.A(\genblk1.pcpi_mul.rs2[0] ),
    .X(_10695_));
 sky130_fd_sc_hd__buf_2 _17393_ (.A(\genblk1.pcpi_mul.rs1[5] ),
    .X(_10696_));
 sky130_fd_sc_hd__buf_2 _17394_ (.A(_10696_),
    .X(_10697_));
 sky130_fd_sc_hd__nand2_1 _17395_ (.A(_10695_),
    .B(_10697_),
    .Y(_10698_));
 sky130_fd_sc_hd__buf_1 _17396_ (.A(\genblk1.pcpi_mul.rs2[4] ),
    .X(_10699_));
 sky130_fd_sc_hd__buf_2 _17397_ (.A(_10699_),
    .X(_10700_));
 sky130_fd_sc_hd__buf_1 _17398_ (.A(\genblk1.pcpi_mul.rs2[5] ),
    .X(_10701_));
 sky130_fd_sc_hd__buf_2 _17399_ (.A(_10701_),
    .X(_10702_));
 sky130_fd_sc_hd__and4_2 _17400_ (.A(_10587_),
    .B(_10594_),
    .C(_10700_),
    .D(_10702_),
    .X(_10703_));
 sky130_fd_sc_hd__clkbuf_2 _17401_ (.A(\genblk1.pcpi_mul.rs1[1] ),
    .X(_10704_));
 sky130_fd_sc_hd__buf_2 _17402_ (.A(_10704_),
    .X(_10705_));
 sky130_fd_sc_hd__buf_1 _17403_ (.A(\genblk1.pcpi_mul.rs2[5] ),
    .X(_10706_));
 sky130_fd_sc_hd__clkbuf_2 _17404_ (.A(_10706_),
    .X(_10707_));
 sky130_fd_sc_hd__buf_2 _17405_ (.A(_10707_),
    .X(_10708_));
 sky130_fd_sc_hd__clkbuf_2 _17406_ (.A(\genblk1.pcpi_mul.rs1[0] ),
    .X(_10709_));
 sky130_fd_sc_hd__buf_2 _17407_ (.A(_10709_),
    .X(_10710_));
 sky130_fd_sc_hd__a22oi_4 _17408_ (.A1(_10705_),
    .A2(_10671_),
    .B1(_10708_),
    .B2(_10710_),
    .Y(_10711_));
 sky130_fd_sc_hd__or3_1 _17409_ (.A(_10698_),
    .B(_10703_),
    .C(_10711_),
    .X(_10712_));
 sky130_fd_sc_hd__o21ai_1 _17410_ (.A1(_10703_),
    .A2(_10711_),
    .B1(_10698_),
    .Y(_10713_));
 sky130_fd_sc_hd__nand3_1 _17411_ (.A(_10673_),
    .B(_10712_),
    .C(_10713_),
    .Y(_10714_));
 sky130_fd_sc_hd__a21o_1 _17412_ (.A1(_10712_),
    .A2(_10713_),
    .B1(_10673_),
    .X(_10715_));
 sky130_fd_sc_hd__nand2_1 _17413_ (.A(_10608_),
    .B(_10644_),
    .Y(_10716_));
 sky130_fd_sc_hd__buf_2 _17414_ (.A(_10647_),
    .X(_10717_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17415_ (.A(\genblk1.pcpi_mul.rs1[4] ),
    .X(_10718_));
 sky130_fd_sc_hd__clkbuf_2 _17416_ (.A(_10718_),
    .X(_10719_));
 sky130_fd_sc_hd__and4_2 _17417_ (.A(_10599_),
    .B(_10631_),
    .C(_10717_),
    .D(_10719_),
    .X(_10720_));
 sky130_fd_sc_hd__clkbuf_4 _17418_ (.A(_10719_),
    .X(_10721_));
 sky130_fd_sc_hd__a22oi_2 _17419_ (.A1(_10611_),
    .A2(_10649_),
    .B1(_10721_),
    .B2(_10640_),
    .Y(_10722_));
 sky130_fd_sc_hd__or2_1 _17420_ (.A(_10720_),
    .B(_10722_),
    .X(_10723_));
 sky130_fd_sc_hd__xor2_1 _17421_ (.A(_10716_),
    .B(_10723_),
    .X(_10724_));
 sky130_fd_sc_hd__nand3_1 _17422_ (.A(_10714_),
    .B(_10715_),
    .C(_10724_),
    .Y(_10725_));
 sky130_fd_sc_hd__a21o_1 _17423_ (.A1(_10714_),
    .A2(_10715_),
    .B1(_10724_),
    .X(_10726_));
 sky130_fd_sc_hd__nand3b_1 _17424_ (.A_N(_10682_),
    .B(_10725_),
    .C(_10726_),
    .Y(_10727_));
 sky130_fd_sc_hd__a21bo_1 _17425_ (.A1(_10725_),
    .A2(_10726_),
    .B1_N(_10682_),
    .X(_10728_));
 sky130_fd_sc_hd__nand3_1 _17426_ (.A(_10694_),
    .B(_10727_),
    .C(_10728_),
    .Y(_10729_));
 sky130_fd_sc_hd__a21o_1 _17427_ (.A1(_10727_),
    .A2(_10728_),
    .B1(_10694_),
    .X(_10730_));
 sky130_fd_sc_hd__and3_1 _17428_ (.A(_10693_),
    .B(_10729_),
    .C(_10730_),
    .X(_10731_));
 sky130_fd_sc_hd__a21o_1 _17429_ (.A1(_10729_),
    .A2(_10730_),
    .B1(_10693_),
    .X(_10732_));
 sky130_fd_sc_hd__and2b_1 _17430_ (.A_N(_10731_),
    .B(_10732_),
    .X(_10733_));
 sky130_fd_sc_hd__and4b_1 _17431_ (.A_N(_10690_),
    .B(_10691_),
    .C(_10733_),
    .D(_10659_),
    .X(_10734_));
 sky130_fd_sc_hd__buf_2 _17432_ (.A(\genblk1.pcpi_mul.rs2[6] ),
    .X(_10735_));
 sky130_fd_sc_hd__clkbuf_4 _17433_ (.A(_10735_),
    .X(_10736_));
 sky130_fd_sc_hd__buf_2 _17434_ (.A(_10736_),
    .X(_10737_));
 sky130_fd_sc_hd__buf_4 _17435_ (.A(_10737_),
    .X(_10738_));
 sky130_fd_sc_hd__nor2_1 _17436_ (.A(_10716_),
    .B(_10723_),
    .Y(_10739_));
 sky130_fd_sc_hd__buf_4 _17437_ (.A(\genblk1.pcpi_mul.rs2[2] ),
    .X(_10740_));
 sky130_fd_sc_hd__buf_2 _17438_ (.A(_10718_),
    .X(_10741_));
 sky130_fd_sc_hd__buf_2 _17439_ (.A(_10741_),
    .X(_10742_));
 sky130_fd_sc_hd__nand4_2 _17440_ (.A(_10640_),
    .B(_10740_),
    .C(_10742_),
    .D(_10697_),
    .Y(_10743_));
 sky130_fd_sc_hd__clkbuf_4 _17441_ (.A(_10664_),
    .X(_10744_));
 sky130_fd_sc_hd__clkbuf_2 _17442_ (.A(\genblk1.pcpi_mul.rs1[5] ),
    .X(_10745_));
 sky130_fd_sc_hd__buf_2 _17443_ (.A(_10745_),
    .X(_10746_));
 sky130_fd_sc_hd__clkbuf_4 _17444_ (.A(_10639_),
    .X(_10747_));
 sky130_fd_sc_hd__a22o_1 _17445_ (.A1(_10631_),
    .A2(_10744_),
    .B1(_10746_),
    .B2(_10747_),
    .X(_10748_));
 sky130_fd_sc_hd__nand2_1 _17446_ (.A(_10743_),
    .B(_10748_),
    .Y(_10749_));
 sky130_fd_sc_hd__nand2_1 _17447_ (.A(_10650_),
    .B(_10644_),
    .Y(_10750_));
 sky130_fd_sc_hd__xor2_1 _17448_ (.A(_10749_),
    .B(_10750_),
    .X(_10751_));
 sky130_fd_sc_hd__buf_1 _17449_ (.A(\genblk1.pcpi_mul.rs1[2] ),
    .X(_10752_));
 sky130_fd_sc_hd__and4_1 _17450_ (.A(_10634_),
    .B(_10752_),
    .C(_10661_),
    .D(_10707_),
    .X(_10753_));
 sky130_fd_sc_hd__buf_2 _17451_ (.A(\genblk1.pcpi_mul.rs1[2] ),
    .X(_10754_));
 sky130_fd_sc_hd__a22oi_2 _17452_ (.A1(_10754_),
    .A2(_10700_),
    .B1(_10702_),
    .B2(_10594_),
    .Y(_10755_));
 sky130_fd_sc_hd__clkbuf_2 _17453_ (.A(\genblk1.pcpi_mul.rs1[6] ),
    .X(_10756_));
 sky130_fd_sc_hd__clkbuf_4 _17454_ (.A(_10756_),
    .X(_10757_));
 sky130_fd_sc_hd__nand2_1 _17455_ (.A(_10695_),
    .B(_10757_),
    .Y(_10758_));
 sky130_fd_sc_hd__or3_2 _17456_ (.A(_10753_),
    .B(_10755_),
    .C(_10758_),
    .X(_10759_));
 sky130_fd_sc_hd__o21ai_2 _17457_ (.A1(_10753_),
    .A2(_10755_),
    .B1(_10758_),
    .Y(_10760_));
 sky130_fd_sc_hd__o21bai_1 _17458_ (.A1(_10698_),
    .A2(_10711_),
    .B1_N(_10703_),
    .Y(_10761_));
 sky130_fd_sc_hd__nand3_1 _17459_ (.A(_10759_),
    .B(_10760_),
    .C(_10761_),
    .Y(_10762_));
 sky130_fd_sc_hd__a21o_1 _17460_ (.A1(_10759_),
    .A2(_10760_),
    .B1(_10761_),
    .X(_10763_));
 sky130_fd_sc_hd__nand3_1 _17461_ (.A(_10751_),
    .B(_10762_),
    .C(_10763_),
    .Y(_10764_));
 sky130_fd_sc_hd__a21o_1 _17462_ (.A1(_10762_),
    .A2(_10763_),
    .B1(_10751_),
    .X(_10765_));
 sky130_fd_sc_hd__a21bo_1 _17463_ (.A1(_10715_),
    .A2(_10724_),
    .B1_N(_10714_),
    .X(_10766_));
 sky130_fd_sc_hd__nand3_2 _17464_ (.A(_10764_),
    .B(_10765_),
    .C(_10766_),
    .Y(_10767_));
 sky130_fd_sc_hd__a21o_1 _17465_ (.A1(_10764_),
    .A2(_10765_),
    .B1(_10766_),
    .X(_10768_));
 sky130_fd_sc_hd__o211ai_2 _17466_ (.A1(_10720_),
    .A2(_10739_),
    .B1(_10767_),
    .C1(_10768_),
    .Y(_10769_));
 sky130_fd_sc_hd__a211o_1 _17467_ (.A1(_10767_),
    .A2(_10768_),
    .B1(_10720_),
    .C1(_10739_),
    .X(_10770_));
 sky130_fd_sc_hd__nand4_2 _17468_ (.A(_10592_),
    .B(_10738_),
    .C(_10769_),
    .D(_10770_),
    .Y(_10771_));
 sky130_fd_sc_hd__a22o_1 _17469_ (.A1(_10592_),
    .A2(_10738_),
    .B1(_10769_),
    .B2(_10770_),
    .X(_10772_));
 sky130_fd_sc_hd__nand2_1 _17470_ (.A(_10727_),
    .B(_10729_),
    .Y(_10773_));
 sky130_fd_sc_hd__nand3_1 _17471_ (.A(_10771_),
    .B(_10772_),
    .C(_10773_),
    .Y(_10774_));
 sky130_fd_sc_hd__a21o_1 _17472_ (.A1(_10771_),
    .A2(_10772_),
    .B1(_10773_),
    .X(_10775_));
 sky130_fd_sc_hd__and2_1 _17473_ (.A(_10774_),
    .B(_10775_),
    .X(_10776_));
 sky130_fd_sc_hd__and3b_1 _17474_ (.A_N(_10731_),
    .B(_10732_),
    .C(_10690_),
    .X(_10777_));
 sky130_fd_sc_hd__nor2_1 _17475_ (.A(_10731_),
    .B(_10777_),
    .Y(_10778_));
 sky130_fd_sc_hd__xnor2_1 _17476_ (.A(_10776_),
    .B(_10778_),
    .Y(_10779_));
 sky130_fd_sc_hd__xor2_1 _17477_ (.A(_10734_),
    .B(_10779_),
    .X(_00110_));
 sky130_fd_sc_hd__a22o_1 _17478_ (.A1(_10777_),
    .A2(_10776_),
    .B1(_10779_),
    .B2(_10734_),
    .X(_10780_));
 sky130_fd_sc_hd__clkbuf_2 _17479_ (.A(\genblk1.pcpi_mul.rs2[7] ),
    .X(_10781_));
 sky130_fd_sc_hd__buf_2 _17480_ (.A(_10781_),
    .X(_10782_));
 sky130_fd_sc_hd__buf_2 _17481_ (.A(_10782_),
    .X(_10783_));
 sky130_fd_sc_hd__buf_4 _17482_ (.A(_10783_),
    .X(_10784_));
 sky130_fd_sc_hd__a22oi_2 _17483_ (.A1(_10598_),
    .A2(_10738_),
    .B1(_10784_),
    .B2(_10591_),
    .Y(_10785_));
 sky130_fd_sc_hd__buf_2 _17484_ (.A(_10704_),
    .X(_10786_));
 sky130_fd_sc_hd__buf_2 _17485_ (.A(\genblk1.pcpi_mul.rs2[6] ),
    .X(_10787_));
 sky130_fd_sc_hd__and4_2 _17486_ (.A(_10587_),
    .B(_10786_),
    .C(_10787_),
    .D(_10782_),
    .X(_10788_));
 sky130_fd_sc_hd__or2_1 _17487_ (.A(_10749_),
    .B(_10750_),
    .X(_10789_));
 sky130_fd_sc_hd__buf_2 _17488_ (.A(_10745_),
    .X(_10790_));
 sky130_fd_sc_hd__nand4_2 _17489_ (.A(_10747_),
    .B(_10631_),
    .C(_10757_),
    .D(_10790_),
    .Y(_10791_));
 sky130_fd_sc_hd__buf_2 _17490_ (.A(_10756_),
    .X(_10792_));
 sky130_fd_sc_hd__clkbuf_2 _17491_ (.A(\genblk1.pcpi_mul.rs1[5] ),
    .X(_10793_));
 sky130_fd_sc_hd__clkbuf_2 _17492_ (.A(_10793_),
    .X(_10794_));
 sky130_fd_sc_hd__a22o_1 _17493_ (.A1(_10599_),
    .A2(_10792_),
    .B1(_10794_),
    .B2(_10610_),
    .X(_10795_));
 sky130_fd_sc_hd__nand2_1 _17494_ (.A(_10791_),
    .B(_10795_),
    .Y(_10796_));
 sky130_fd_sc_hd__buf_2 _17495_ (.A(_10665_),
    .X(_10797_));
 sky130_fd_sc_hd__nand2_1 _17496_ (.A(_10624_),
    .B(_10797_),
    .Y(_10798_));
 sky130_fd_sc_hd__xor2_1 _17497_ (.A(_10796_),
    .B(_10798_),
    .X(_10799_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17498_ (.A(\genblk1.pcpi_mul.rs1[3] ),
    .X(_10800_));
 sky130_fd_sc_hd__and4_1 _17499_ (.A(_10752_),
    .B(_10800_),
    .C(_10670_),
    .D(_10701_),
    .X(_10801_));
 sky130_fd_sc_hd__buf_2 _17500_ (.A(\genblk1.pcpi_mul.rs2[4] ),
    .X(_10802_));
 sky130_fd_sc_hd__buf_2 _17501_ (.A(_10706_),
    .X(_10803_));
 sky130_fd_sc_hd__a22oi_2 _17502_ (.A1(_10648_),
    .A2(_10802_),
    .B1(_10803_),
    .B2(_10628_),
    .Y(_10804_));
 sky130_fd_sc_hd__buf_2 _17503_ (.A(\genblk1.pcpi_mul.rs1[7] ),
    .X(_10805_));
 sky130_fd_sc_hd__nand2_1 _17504_ (.A(_10582_),
    .B(_10805_),
    .Y(_10806_));
 sky130_fd_sc_hd__or3_1 _17505_ (.A(_10801_),
    .B(_10804_),
    .C(_10806_),
    .X(_10807_));
 sky130_fd_sc_hd__o21ai_1 _17506_ (.A1(_10801_),
    .A2(_10804_),
    .B1(_10806_),
    .Y(_10808_));
 sky130_fd_sc_hd__o21bai_1 _17507_ (.A1(_10755_),
    .A2(_10758_),
    .B1_N(_10753_),
    .Y(_10809_));
 sky130_fd_sc_hd__nand3_1 _17508_ (.A(_10807_),
    .B(_10808_),
    .C(_10809_),
    .Y(_10810_));
 sky130_fd_sc_hd__a21o_1 _17509_ (.A1(_10807_),
    .A2(_10808_),
    .B1(_10809_),
    .X(_10811_));
 sky130_fd_sc_hd__nand3_2 _17510_ (.A(_10799_),
    .B(_10810_),
    .C(_10811_),
    .Y(_10812_));
 sky130_fd_sc_hd__a21o_1 _17511_ (.A1(_10810_),
    .A2(_10811_),
    .B1(_10799_),
    .X(_10813_));
 sky130_fd_sc_hd__a21bo_1 _17512_ (.A1(_10751_),
    .A2(_10763_),
    .B1_N(_10762_),
    .X(_10814_));
 sky130_fd_sc_hd__and3_1 _17513_ (.A(_10812_),
    .B(_10813_),
    .C(_10814_),
    .X(_10815_));
 sky130_fd_sc_hd__a21oi_1 _17514_ (.A1(_10812_),
    .A2(_10813_),
    .B1(_10814_),
    .Y(_10816_));
 sky130_fd_sc_hd__a211oi_2 _17515_ (.A1(_10743_),
    .A2(_10789_),
    .B1(_10815_),
    .C1(_10816_),
    .Y(_10817_));
 sky130_fd_sc_hd__o211a_1 _17516_ (.A1(_10815_),
    .A2(_10816_),
    .B1(_10743_),
    .C1(_10789_),
    .X(_10818_));
 sky130_fd_sc_hd__nor4_2 _17517_ (.A(_10785_),
    .B(_10788_),
    .C(_10817_),
    .D(_10818_),
    .Y(_10819_));
 sky130_fd_sc_hd__o22a_1 _17518_ (.A1(_10785_),
    .A2(_10788_),
    .B1(_10817_),
    .B2(_10818_),
    .X(_10820_));
 sky130_fd_sc_hd__or3_2 _17519_ (.A(_10771_),
    .B(_10819_),
    .C(_10820_),
    .X(_10821_));
 sky130_fd_sc_hd__o21ai_1 _17520_ (.A1(_10819_),
    .A2(_10820_),
    .B1(_10771_),
    .Y(_10822_));
 sky130_fd_sc_hd__nand2_1 _17521_ (.A(_10767_),
    .B(_10769_),
    .Y(_10823_));
 sky130_fd_sc_hd__and3_1 _17522_ (.A(_10821_),
    .B(_10822_),
    .C(_10823_),
    .X(_10824_));
 sky130_fd_sc_hd__a21oi_1 _17523_ (.A1(_10821_),
    .A2(_10822_),
    .B1(_10823_),
    .Y(_10825_));
 sky130_fd_sc_hd__nor2_1 _17524_ (.A(_10824_),
    .B(_10825_),
    .Y(_10826_));
 sky130_vsdinv _17525_ (.A(_10774_),
    .Y(_10827_));
 sky130_fd_sc_hd__and3_1 _17526_ (.A(_10731_),
    .B(_10774_),
    .C(_10775_),
    .X(_10828_));
 sky130_fd_sc_hd__nor2_1 _17527_ (.A(_10827_),
    .B(_10828_),
    .Y(_10829_));
 sky130_fd_sc_hd__xnor2_1 _17528_ (.A(_10826_),
    .B(_10829_),
    .Y(_10830_));
 sky130_fd_sc_hd__nand2_1 _17529_ (.A(_10780_),
    .B(_10830_),
    .Y(_10831_));
 sky130_fd_sc_hd__or2_1 _17530_ (.A(_10780_),
    .B(_10830_),
    .X(_10832_));
 sky130_fd_sc_hd__and2_1 _17531_ (.A(_10831_),
    .B(_10832_),
    .X(_10833_));
 sky130_fd_sc_hd__clkbuf_1 _17532_ (.A(_10833_),
    .X(_00111_));
 sky130_fd_sc_hd__nand2_1 _17533_ (.A(_10826_),
    .B(_10828_),
    .Y(_10834_));
 sky130_fd_sc_hd__nand2_1 _17534_ (.A(_10827_),
    .B(_10826_),
    .Y(_10835_));
 sky130_fd_sc_hd__clkbuf_4 _17535_ (.A(\genblk1.pcpi_mul.rs2[7] ),
    .X(_10836_));
 sky130_fd_sc_hd__buf_2 _17536_ (.A(\genblk1.pcpi_mul.rs2[8] ),
    .X(_10837_));
 sky130_fd_sc_hd__nand4_2 _17537_ (.A(_10709_),
    .B(_10704_),
    .C(_10836_),
    .D(_10837_),
    .Y(_10838_));
 sky130_fd_sc_hd__clkbuf_4 _17538_ (.A(\genblk1.pcpi_mul.rs2[8] ),
    .X(_10839_));
 sky130_fd_sc_hd__a22o_1 _17539_ (.A1(\genblk1.pcpi_mul.rs1[1] ),
    .A2(_10781_),
    .B1(_10839_),
    .B2(\genblk1.pcpi_mul.rs1[0] ),
    .X(_10840_));
 sky130_fd_sc_hd__and2_1 _17540_ (.A(_10606_),
    .B(\genblk1.pcpi_mul.rs2[6] ),
    .X(_10841_));
 sky130_fd_sc_hd__nand3_1 _17541_ (.A(_10838_),
    .B(_10840_),
    .C(_10841_),
    .Y(_10842_));
 sky130_fd_sc_hd__a21o_1 _17542_ (.A1(_10838_),
    .A2(_10840_),
    .B1(_10841_),
    .X(_10843_));
 sky130_fd_sc_hd__and3_1 _17543_ (.A(_10788_),
    .B(_10842_),
    .C(_10843_),
    .X(_10844_));
 sky130_fd_sc_hd__a21oi_1 _17544_ (.A1(_10842_),
    .A2(_10843_),
    .B1(_10788_),
    .Y(_10845_));
 sky130_fd_sc_hd__or2_1 _17545_ (.A(_10844_),
    .B(_10845_),
    .X(_10846_));
 sky130_fd_sc_hd__or2_1 _17546_ (.A(_10796_),
    .B(_10798_),
    .X(_10847_));
 sky130_fd_sc_hd__clkbuf_4 _17547_ (.A(\genblk1.pcpi_mul.rs1[6] ),
    .X(_10848_));
 sky130_fd_sc_hd__clkbuf_2 _17548_ (.A(\genblk1.pcpi_mul.rs1[7] ),
    .X(_10849_));
 sky130_fd_sc_hd__and4_2 _17549_ (.A(\genblk1.pcpi_mul.rs2[1] ),
    .B(\genblk1.pcpi_mul.rs2[2] ),
    .C(_10848_),
    .D(_10849_),
    .X(_10850_));
 sky130_fd_sc_hd__clkbuf_2 _17550_ (.A(\genblk1.pcpi_mul.rs1[7] ),
    .X(_10851_));
 sky130_fd_sc_hd__buf_2 _17551_ (.A(_10851_),
    .X(_10852_));
 sky130_fd_sc_hd__a22oi_1 _17552_ (.A1(_10610_),
    .A2(_10792_),
    .B1(_10852_),
    .B2(_10599_),
    .Y(_10853_));
 sky130_fd_sc_hd__or2_1 _17553_ (.A(_10850_),
    .B(_10853_),
    .X(_10854_));
 sky130_fd_sc_hd__buf_2 _17554_ (.A(_10794_),
    .X(_10855_));
 sky130_fd_sc_hd__nand2_1 _17555_ (.A(_10624_),
    .B(_10855_),
    .Y(_10856_));
 sky130_fd_sc_hd__xor2_1 _17556_ (.A(_10854_),
    .B(_10856_),
    .X(_10857_));
 sky130_fd_sc_hd__buf_2 _17557_ (.A(\genblk1.pcpi_mul.rs1[8] ),
    .X(_10858_));
 sky130_fd_sc_hd__nand2_1 _17558_ (.A(_10582_),
    .B(_10858_),
    .Y(_10859_));
 sky130_fd_sc_hd__and4_1 _17559_ (.A(_10800_),
    .B(_10670_),
    .C(_10664_),
    .D(_10701_),
    .X(_10860_));
 sky130_fd_sc_hd__clkbuf_2 _17560_ (.A(_10647_),
    .X(_10861_));
 sky130_fd_sc_hd__a22oi_2 _17561_ (.A1(_10661_),
    .A2(_10741_),
    .B1(_10803_),
    .B2(_10861_),
    .Y(_10862_));
 sky130_fd_sc_hd__or3_1 _17562_ (.A(_10859_),
    .B(_10860_),
    .C(_10862_),
    .X(_10863_));
 sky130_fd_sc_hd__o21ai_1 _17563_ (.A1(_10860_),
    .A2(_10862_),
    .B1(_10859_),
    .Y(_10864_));
 sky130_fd_sc_hd__o21bai_1 _17564_ (.A1(_10804_),
    .A2(_10806_),
    .B1_N(_10801_),
    .Y(_10865_));
 sky130_fd_sc_hd__nand3_1 _17565_ (.A(_10863_),
    .B(_10864_),
    .C(_10865_),
    .Y(_10866_));
 sky130_fd_sc_hd__a21o_1 _17566_ (.A1(_10863_),
    .A2(_10864_),
    .B1(_10865_),
    .X(_10867_));
 sky130_fd_sc_hd__nand3_1 _17567_ (.A(_10857_),
    .B(_10866_),
    .C(_10867_),
    .Y(_10868_));
 sky130_fd_sc_hd__a21o_1 _17568_ (.A1(_10866_),
    .A2(_10867_),
    .B1(_10857_),
    .X(_10869_));
 sky130_fd_sc_hd__a21bo_1 _17569_ (.A1(_10799_),
    .A2(_10811_),
    .B1_N(_10810_),
    .X(_10870_));
 sky130_fd_sc_hd__and3_1 _17570_ (.A(_10868_),
    .B(_10869_),
    .C(_10870_),
    .X(_10871_));
 sky130_fd_sc_hd__a21oi_1 _17571_ (.A1(_10868_),
    .A2(_10869_),
    .B1(_10870_),
    .Y(_10872_));
 sky130_fd_sc_hd__a211oi_2 _17572_ (.A1(_10791_),
    .A2(_10847_),
    .B1(_10871_),
    .C1(_10872_),
    .Y(_10873_));
 sky130_fd_sc_hd__o211a_1 _17573_ (.A1(_10871_),
    .A2(_10872_),
    .B1(_10791_),
    .C1(_10847_),
    .X(_10874_));
 sky130_fd_sc_hd__or3_2 _17574_ (.A(_10846_),
    .B(_10873_),
    .C(_10874_),
    .X(_10875_));
 sky130_fd_sc_hd__o21ai_2 _17575_ (.A1(_10873_),
    .A2(_10874_),
    .B1(_10846_),
    .Y(_10876_));
 sky130_fd_sc_hd__and3_1 _17576_ (.A(_10819_),
    .B(_10875_),
    .C(_10876_),
    .X(_10877_));
 sky130_fd_sc_hd__a21oi_1 _17577_ (.A1(_10875_),
    .A2(_10876_),
    .B1(_10819_),
    .Y(_10878_));
 sky130_fd_sc_hd__or2_1 _17578_ (.A(_10877_),
    .B(_10878_),
    .X(_10879_));
 sky130_fd_sc_hd__nor2_1 _17579_ (.A(_10815_),
    .B(_10817_),
    .Y(_10880_));
 sky130_fd_sc_hd__xnor2_1 _17580_ (.A(_10821_),
    .B(_10880_),
    .Y(_10881_));
 sky130_fd_sc_hd__xnor2_1 _17581_ (.A(_10879_),
    .B(_10881_),
    .Y(_10882_));
 sky130_fd_sc_hd__xor2_1 _17582_ (.A(_10824_),
    .B(_10882_),
    .X(_10883_));
 sky130_fd_sc_hd__xor2_1 _17583_ (.A(_10835_),
    .B(_10883_),
    .X(_10884_));
 sky130_fd_sc_hd__a21bo_1 _17584_ (.A1(_10834_),
    .A2(_10831_),
    .B1_N(_10884_),
    .X(_10885_));
 sky130_fd_sc_hd__a221o_1 _17585_ (.A1(_10826_),
    .A2(_10828_),
    .B1(_10830_),
    .B2(_10780_),
    .C1(_10884_),
    .X(_10886_));
 sky130_fd_sc_hd__and2_1 _17586_ (.A(_10885_),
    .B(_10886_),
    .X(_10887_));
 sky130_fd_sc_hd__clkbuf_1 _17587_ (.A(_10887_),
    .X(_00112_));
 sky130_fd_sc_hd__nor2_1 _17588_ (.A(_10835_),
    .B(_10883_),
    .Y(_10888_));
 sky130_vsdinv _17589_ (.A(_10888_),
    .Y(_10889_));
 sky130_fd_sc_hd__and4b_1 _17590_ (.A_N(_10882_),
    .B(_10823_),
    .C(_10822_),
    .D(_10821_),
    .X(_10890_));
 sky130_fd_sc_hd__or2_1 _17591_ (.A(_10821_),
    .B(_10880_),
    .X(_10891_));
 sky130_fd_sc_hd__clkbuf_2 _17592_ (.A(\genblk1.pcpi_mul.rs2[9] ),
    .X(_10892_));
 sky130_fd_sc_hd__clkbuf_4 _17593_ (.A(_10892_),
    .X(_10893_));
 sky130_fd_sc_hd__clkbuf_2 _17594_ (.A(_10893_),
    .X(_10894_));
 sky130_fd_sc_hd__buf_4 _17595_ (.A(_10894_),
    .X(_10895_));
 sky130_fd_sc_hd__and4_1 _17596_ (.A(\genblk1.pcpi_mul.rs1[1] ),
    .B(\genblk1.pcpi_mul.rs1[2] ),
    .C(_10781_),
    .D(\genblk1.pcpi_mul.rs2[8] ),
    .X(_10896_));
 sky130_fd_sc_hd__a22oi_2 _17597_ (.A1(_10606_),
    .A2(_10836_),
    .B1(_10837_),
    .B2(_10704_),
    .Y(_10897_));
 sky130_fd_sc_hd__and4bb_1 _17598_ (.A_N(_10896_),
    .B_N(_10897_),
    .C(_10861_),
    .D(_10735_),
    .X(_10898_));
 sky130_fd_sc_hd__o2bb2a_1 _17599_ (.A1_N(_10861_),
    .A2_N(_10735_),
    .B1(_10896_),
    .B2(_10897_),
    .X(_10899_));
 sky130_fd_sc_hd__a21bo_1 _17600_ (.A1(_10840_),
    .A2(_10841_),
    .B1_N(_10838_),
    .X(_10900_));
 sky130_fd_sc_hd__or3b_2 _17601_ (.A(_10898_),
    .B(_10899_),
    .C_N(_10900_),
    .X(_10901_));
 sky130_fd_sc_hd__o21bai_1 _17602_ (.A1(_10898_),
    .A2(_10899_),
    .B1_N(_10900_),
    .Y(_10902_));
 sky130_fd_sc_hd__and3_1 _17603_ (.A(_10844_),
    .B(_10901_),
    .C(_10902_),
    .X(_10903_));
 sky130_vsdinv _17604_ (.A(_10903_),
    .Y(_10904_));
 sky130_fd_sc_hd__a21o_1 _17605_ (.A1(_10901_),
    .A2(_10902_),
    .B1(_10844_),
    .X(_10905_));
 sky130_fd_sc_hd__nor2_1 _17606_ (.A(_10854_),
    .B(_10856_),
    .Y(_10906_));
 sky130_fd_sc_hd__buf_2 _17607_ (.A(\genblk1.pcpi_mul.rs1[8] ),
    .X(_10907_));
 sky130_fd_sc_hd__and4_1 _17608_ (.A(\genblk1.pcpi_mul.rs2[1] ),
    .B(\genblk1.pcpi_mul.rs2[2] ),
    .C(_10849_),
    .D(_10907_),
    .X(_10908_));
 sky130_fd_sc_hd__buf_2 _17609_ (.A(\genblk1.pcpi_mul.rs1[7] ),
    .X(_10909_));
 sky130_fd_sc_hd__a22oi_1 _17610_ (.A1(\genblk1.pcpi_mul.rs2[2] ),
    .A2(_10909_),
    .B1(_10858_),
    .B2(_10639_),
    .Y(_10910_));
 sky130_fd_sc_hd__or2_1 _17611_ (.A(_10908_),
    .B(_10910_),
    .X(_10911_));
 sky130_fd_sc_hd__buf_2 _17612_ (.A(_10792_),
    .X(_10912_));
 sky130_fd_sc_hd__nand2_1 _17613_ (.A(_10624_),
    .B(_10912_),
    .Y(_10913_));
 sky130_fd_sc_hd__xor2_1 _17614_ (.A(_10911_),
    .B(_10913_),
    .X(_10914_));
 sky130_fd_sc_hd__and4_1 _17615_ (.A(_10699_),
    .B(_10664_),
    .C(_10701_),
    .D(_10793_),
    .X(_10915_));
 sky130_fd_sc_hd__buf_2 _17616_ (.A(_10706_),
    .X(_10916_));
 sky130_fd_sc_hd__a22oi_2 _17617_ (.A1(_10741_),
    .A2(_10916_),
    .B1(_10696_),
    .B2(_10802_),
    .Y(_10917_));
 sky130_fd_sc_hd__clkbuf_2 _17618_ (.A(\genblk1.pcpi_mul.rs1[9] ),
    .X(_10918_));
 sky130_fd_sc_hd__buf_2 _17619_ (.A(_10918_),
    .X(_10919_));
 sky130_fd_sc_hd__nand2_1 _17620_ (.A(_10582_),
    .B(_10919_),
    .Y(_10920_));
 sky130_fd_sc_hd__or3_1 _17621_ (.A(_10915_),
    .B(_10917_),
    .C(_10920_),
    .X(_10921_));
 sky130_fd_sc_hd__o21ai_1 _17622_ (.A1(_10915_),
    .A2(_10917_),
    .B1(_10920_),
    .Y(_10922_));
 sky130_fd_sc_hd__o21bai_1 _17623_ (.A1(_10859_),
    .A2(_10862_),
    .B1_N(_10860_),
    .Y(_10923_));
 sky130_fd_sc_hd__nand3_1 _17624_ (.A(_10921_),
    .B(_10922_),
    .C(_10923_),
    .Y(_10924_));
 sky130_fd_sc_hd__a21o_1 _17625_ (.A1(_10921_),
    .A2(_10922_),
    .B1(_10923_),
    .X(_10925_));
 sky130_fd_sc_hd__nand3_1 _17626_ (.A(_10914_),
    .B(_10924_),
    .C(_10925_),
    .Y(_10926_));
 sky130_fd_sc_hd__a21o_1 _17627_ (.A1(_10924_),
    .A2(_10925_),
    .B1(_10914_),
    .X(_10927_));
 sky130_fd_sc_hd__a21bo_1 _17628_ (.A1(_10857_),
    .A2(_10867_),
    .B1_N(_10866_),
    .X(_10928_));
 sky130_fd_sc_hd__nand3_2 _17629_ (.A(_10926_),
    .B(_10927_),
    .C(_10928_),
    .Y(_10929_));
 sky130_fd_sc_hd__a21o_1 _17630_ (.A1(_10926_),
    .A2(_10927_),
    .B1(_10928_),
    .X(_10930_));
 sky130_fd_sc_hd__o211ai_4 _17631_ (.A1(_10850_),
    .A2(_10906_),
    .B1(_10929_),
    .C1(_10930_),
    .Y(_10931_));
 sky130_fd_sc_hd__a211o_1 _17632_ (.A1(_10929_),
    .A2(_10930_),
    .B1(_10850_),
    .C1(_10906_),
    .X(_10932_));
 sky130_fd_sc_hd__and4_2 _17633_ (.A(_10904_),
    .B(_10905_),
    .C(_10931_),
    .D(_10932_),
    .X(_10933_));
 sky130_fd_sc_hd__a22oi_4 _17634_ (.A1(_10904_),
    .A2(_10905_),
    .B1(_10931_),
    .B2(_10932_),
    .Y(_10934_));
 sky130_fd_sc_hd__or3_2 _17635_ (.A(_10875_),
    .B(_10933_),
    .C(_10934_),
    .X(_10935_));
 sky130_fd_sc_hd__o21ai_1 _17636_ (.A1(_10933_),
    .A2(_10934_),
    .B1(_10875_),
    .Y(_10936_));
 sky130_fd_sc_hd__nand4_1 _17637_ (.A(_10603_),
    .B(_10895_),
    .C(_10935_),
    .D(_10936_),
    .Y(_10937_));
 sky130_fd_sc_hd__a22o_1 _17638_ (.A1(_10603_),
    .A2(_10895_),
    .B1(_10935_),
    .B2(_10936_),
    .X(_10938_));
 sky130_fd_sc_hd__nor2_2 _17639_ (.A(_10871_),
    .B(_10873_),
    .Y(_10939_));
 sky130_fd_sc_hd__xnor2_1 _17640_ (.A(_10877_),
    .B(_10939_),
    .Y(_10940_));
 sky130_fd_sc_hd__and3_1 _17641_ (.A(_10937_),
    .B(_10938_),
    .C(_10940_),
    .X(_10941_));
 sky130_fd_sc_hd__a21oi_1 _17642_ (.A1(_10937_),
    .A2(_10938_),
    .B1(_10940_),
    .Y(_10942_));
 sky130_fd_sc_hd__or2_1 _17643_ (.A(_10941_),
    .B(_10942_),
    .X(_10943_));
 sky130_fd_sc_hd__or2_1 _17644_ (.A(_10891_),
    .B(_10943_),
    .X(_10944_));
 sky130_fd_sc_hd__or2_1 _17645_ (.A(_10879_),
    .B(_10881_),
    .X(_10945_));
 sky130_fd_sc_hd__or3_1 _17646_ (.A(_10945_),
    .B(_10941_),
    .C(_10942_),
    .X(_10946_));
 sky130_fd_sc_hd__o21ai_1 _17647_ (.A1(_10941_),
    .A2(_10942_),
    .B1(_10945_),
    .Y(_10947_));
 sky130_fd_sc_hd__a21bo_1 _17648_ (.A1(_10946_),
    .A2(_10947_),
    .B1_N(_10891_),
    .X(_10948_));
 sky130_fd_sc_hd__and3_1 _17649_ (.A(_10890_),
    .B(_10944_),
    .C(_10948_),
    .X(_10949_));
 sky130_fd_sc_hd__a21oi_1 _17650_ (.A1(_10944_),
    .A2(_10948_),
    .B1(_10890_),
    .Y(_10950_));
 sky130_fd_sc_hd__a211o_1 _17651_ (.A1(_10889_),
    .A2(_10885_),
    .B1(_10949_),
    .C1(_10950_),
    .X(_10951_));
 sky130_fd_sc_hd__o211ai_1 _17652_ (.A1(_10949_),
    .A2(_10950_),
    .B1(_10889_),
    .C1(_10885_),
    .Y(_10952_));
 sky130_fd_sc_hd__and2_1 _17653_ (.A(_10951_),
    .B(_10952_),
    .X(_10953_));
 sky130_fd_sc_hd__clkbuf_1 _17654_ (.A(_10953_),
    .X(_00113_));
 sky130_vsdinv _17655_ (.A(_10949_),
    .Y(_10954_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17656_ (.A(\genblk1.pcpi_mul.rs2[10] ),
    .X(_10955_));
 sky130_fd_sc_hd__clkbuf_2 _17657_ (.A(_10955_),
    .X(_10956_));
 sky130_fd_sc_hd__clkbuf_4 _17658_ (.A(_10956_),
    .X(_10957_));
 sky130_fd_sc_hd__buf_4 _17659_ (.A(_10957_),
    .X(_10958_));
 sky130_fd_sc_hd__a22oi_2 _17660_ (.A1(_10598_),
    .A2(_10895_),
    .B1(_10958_),
    .B2(_10592_),
    .Y(_10959_));
 sky130_fd_sc_hd__buf_2 _17661_ (.A(\genblk1.pcpi_mul.rs2[9] ),
    .X(_10960_));
 sky130_fd_sc_hd__clkbuf_4 _17662_ (.A(_10960_),
    .X(_10961_));
 sky130_fd_sc_hd__clkbuf_2 _17663_ (.A(\genblk1.pcpi_mul.rs2[10] ),
    .X(_10962_));
 sky130_fd_sc_hd__buf_2 _17664_ (.A(_10962_),
    .X(_10963_));
 sky130_fd_sc_hd__and3_1 _17665_ (.A(_10710_),
    .B(_10705_),
    .C(_10963_),
    .X(_10964_));
 sky130_fd_sc_hd__and2_2 _17666_ (.A(_10961_),
    .B(_10964_),
    .X(_10965_));
 sky130_fd_sc_hd__nor2_1 _17667_ (.A(_10911_),
    .B(_10913_),
    .Y(_10966_));
 sky130_fd_sc_hd__clkbuf_4 _17668_ (.A(_10907_),
    .X(_10967_));
 sky130_fd_sc_hd__clkbuf_2 _17669_ (.A(\genblk1.pcpi_mul.rs1[9] ),
    .X(_10968_));
 sky130_fd_sc_hd__clkbuf_4 _17670_ (.A(_10968_),
    .X(_10969_));
 sky130_fd_sc_hd__nand4_4 _17671_ (.A(_10599_),
    .B(_10631_),
    .C(_10967_),
    .D(_10969_),
    .Y(_10970_));
 sky130_fd_sc_hd__a22o_1 _17672_ (.A1(_10610_),
    .A2(_10858_),
    .B1(_10919_),
    .B2(_10639_),
    .X(_10971_));
 sky130_fd_sc_hd__nand2_1 _17673_ (.A(_10970_),
    .B(_10971_),
    .Y(_10972_));
 sky130_fd_sc_hd__clkbuf_4 _17674_ (.A(_10805_),
    .X(_10973_));
 sky130_fd_sc_hd__nand2_1 _17675_ (.A(_10624_),
    .B(_10973_),
    .Y(_10974_));
 sky130_fd_sc_hd__xor2_1 _17676_ (.A(_10972_),
    .B(_10974_),
    .X(_10975_));
 sky130_fd_sc_hd__clkbuf_2 _17677_ (.A(\genblk1.pcpi_mul.rs1[10] ),
    .X(_10976_));
 sky130_fd_sc_hd__nand2_1 _17678_ (.A(\genblk1.pcpi_mul.rs2[0] ),
    .B(_10976_),
    .Y(_10977_));
 sky130_fd_sc_hd__buf_2 _17679_ (.A(\genblk1.pcpi_mul.rs1[6] ),
    .X(_10978_));
 sky130_fd_sc_hd__and4_1 _17680_ (.A(_10699_),
    .B(_10706_),
    .C(_10978_),
    .D(_10793_),
    .X(_10979_));
 sky130_fd_sc_hd__a22oi_4 _17681_ (.A1(_10670_),
    .A2(_10848_),
    .B1(_10745_),
    .B2(_10916_),
    .Y(_10980_));
 sky130_fd_sc_hd__or3_1 _17682_ (.A(_10977_),
    .B(_10979_),
    .C(_10980_),
    .X(_10981_));
 sky130_fd_sc_hd__o21ai_1 _17683_ (.A1(_10979_),
    .A2(_10980_),
    .B1(_10977_),
    .Y(_10982_));
 sky130_fd_sc_hd__o21bai_1 _17684_ (.A1(_10917_),
    .A2(_10920_),
    .B1_N(_10915_),
    .Y(_10983_));
 sky130_fd_sc_hd__nand3_1 _17685_ (.A(_10981_),
    .B(_10982_),
    .C(_10983_),
    .Y(_10984_));
 sky130_fd_sc_hd__a21o_1 _17686_ (.A1(_10981_),
    .A2(_10982_),
    .B1(_10983_),
    .X(_10985_));
 sky130_fd_sc_hd__nand3_1 _17687_ (.A(_10975_),
    .B(_10984_),
    .C(_10985_),
    .Y(_10986_));
 sky130_fd_sc_hd__a21o_1 _17688_ (.A1(_10984_),
    .A2(_10985_),
    .B1(_10975_),
    .X(_10987_));
 sky130_fd_sc_hd__a21bo_1 _17689_ (.A1(_10914_),
    .A2(_10925_),
    .B1_N(_10924_),
    .X(_10988_));
 sky130_fd_sc_hd__nand3_1 _17690_ (.A(_10986_),
    .B(_10987_),
    .C(_10988_),
    .Y(_10989_));
 sky130_fd_sc_hd__a21o_1 _17691_ (.A1(_10986_),
    .A2(_10987_),
    .B1(_10988_),
    .X(_10990_));
 sky130_fd_sc_hd__o211a_1 _17692_ (.A1(_10908_),
    .A2(_10966_),
    .B1(_10989_),
    .C1(_10990_),
    .X(_10991_));
 sky130_fd_sc_hd__a211oi_2 _17693_ (.A1(_10989_),
    .A2(_10990_),
    .B1(_10908_),
    .C1(_10966_),
    .Y(_10992_));
 sky130_fd_sc_hd__buf_2 _17694_ (.A(_10735_),
    .X(_10993_));
 sky130_fd_sc_hd__nand2_1 _17695_ (.A(_10721_),
    .B(_10993_),
    .Y(_10994_));
 sky130_fd_sc_hd__buf_2 _17696_ (.A(\genblk1.pcpi_mul.rs2[7] ),
    .X(_10995_));
 sky130_fd_sc_hd__and4_1 _17697_ (.A(_10752_),
    .B(_10648_),
    .C(_10995_),
    .D(_10837_),
    .X(_10996_));
 sky130_fd_sc_hd__clkbuf_4 _17698_ (.A(_10781_),
    .X(_10997_));
 sky130_fd_sc_hd__buf_2 _17699_ (.A(_10839_),
    .X(_10998_));
 sky130_fd_sc_hd__a22oi_1 _17700_ (.A1(_10717_),
    .A2(_10997_),
    .B1(_10998_),
    .B2(_10754_),
    .Y(_10999_));
 sky130_fd_sc_hd__nor2_1 _17701_ (.A(_10996_),
    .B(_10999_),
    .Y(_11000_));
 sky130_fd_sc_hd__xnor2_2 _17702_ (.A(_10994_),
    .B(_11000_),
    .Y(_11001_));
 sky130_fd_sc_hd__or2_2 _17703_ (.A(_10896_),
    .B(_10898_),
    .X(_11002_));
 sky130_fd_sc_hd__xnor2_1 _17704_ (.A(_11001_),
    .B(_11002_),
    .Y(_11003_));
 sky130_vsdinv _17705_ (.A(_10901_),
    .Y(_11004_));
 sky130_fd_sc_hd__xor2_1 _17706_ (.A(_11001_),
    .B(_11002_),
    .X(_11005_));
 sky130_fd_sc_hd__or3_1 _17707_ (.A(_11004_),
    .B(_10903_),
    .C(_11005_),
    .X(_11006_));
 sky130_fd_sc_hd__nand2_1 _17708_ (.A(_10903_),
    .B(_11005_),
    .Y(_11007_));
 sky130_fd_sc_hd__o211ai_1 _17709_ (.A1(_10901_),
    .A2(_11003_),
    .B1(_11006_),
    .C1(_11007_),
    .Y(_11008_));
 sky130_fd_sc_hd__or3_2 _17710_ (.A(_10991_),
    .B(_10992_),
    .C(_11008_),
    .X(_11009_));
 sky130_fd_sc_hd__o21ai_1 _17711_ (.A1(_10991_),
    .A2(_10992_),
    .B1(_11008_),
    .Y(_11010_));
 sky130_fd_sc_hd__and3_1 _17712_ (.A(_10933_),
    .B(_11009_),
    .C(_11010_),
    .X(_11011_));
 sky130_fd_sc_hd__a21oi_1 _17713_ (.A1(_11009_),
    .A2(_11010_),
    .B1(_10933_),
    .Y(_11012_));
 sky130_fd_sc_hd__or4_2 _17714_ (.A(_10959_),
    .B(_10965_),
    .C(_11011_),
    .D(_11012_),
    .X(_11013_));
 sky130_fd_sc_hd__o22ai_2 _17715_ (.A1(_10959_),
    .A2(_10965_),
    .B1(_11011_),
    .B2(_11012_),
    .Y(_11014_));
 sky130_fd_sc_hd__nand3b_1 _17716_ (.A_N(_10937_),
    .B(_11013_),
    .C(_11014_),
    .Y(_11015_));
 sky130_fd_sc_hd__a21bo_1 _17717_ (.A1(_11013_),
    .A2(_11014_),
    .B1_N(_10937_),
    .X(_11016_));
 sky130_fd_sc_hd__nand2_2 _17718_ (.A(_10929_),
    .B(_10931_),
    .Y(_11017_));
 sky130_fd_sc_hd__xnor2_1 _17719_ (.A(_10935_),
    .B(_11017_),
    .Y(_11018_));
 sky130_fd_sc_hd__and3_1 _17720_ (.A(_11015_),
    .B(_11016_),
    .C(_11018_),
    .X(_11019_));
 sky130_fd_sc_hd__a21oi_1 _17721_ (.A1(_11015_),
    .A2(_11016_),
    .B1(_11018_),
    .Y(_11020_));
 sky130_fd_sc_hd__o21bai_1 _17722_ (.A1(_11019_),
    .A2(_11020_),
    .B1_N(_10941_),
    .Y(_11021_));
 sky130_fd_sc_hd__or3b_2 _17723_ (.A(_11019_),
    .B(_11020_),
    .C_N(_10941_),
    .X(_11022_));
 sky130_fd_sc_hd__or2b_1 _17724_ (.A(_10939_),
    .B_N(_10877_),
    .X(_11023_));
 sky130_fd_sc_hd__a21bo_1 _17725_ (.A1(_11021_),
    .A2(_11022_),
    .B1_N(_11023_),
    .X(_11024_));
 sky130_fd_sc_hd__nand3b_2 _17726_ (.A_N(_11023_),
    .B(_11021_),
    .C(_11022_),
    .Y(_11025_));
 sky130_fd_sc_hd__a21oi_1 _17727_ (.A1(_10891_),
    .A2(_10945_),
    .B1(_10943_),
    .Y(_11026_));
 sky130_fd_sc_hd__and3_1 _17728_ (.A(_11024_),
    .B(_11025_),
    .C(_11026_),
    .X(_11027_));
 sky130_fd_sc_hd__a21oi_1 _17729_ (.A1(_11024_),
    .A2(_11025_),
    .B1(_11026_),
    .Y(_11028_));
 sky130_fd_sc_hd__a211oi_1 _17730_ (.A1(_10954_),
    .A2(_10951_),
    .B1(_11027_),
    .C1(_11028_),
    .Y(_11029_));
 sky130_fd_sc_hd__o211a_1 _17731_ (.A1(_11027_),
    .A2(_11028_),
    .B1(_10954_),
    .C1(_10951_),
    .X(_11030_));
 sky130_fd_sc_hd__nor2_1 _17732_ (.A(_11029_),
    .B(_11030_),
    .Y(_00056_));
 sky130_fd_sc_hd__or2b_1 _17733_ (.A(_10935_),
    .B_N(_11017_),
    .X(_11031_));
 sky130_vsdinv _17734_ (.A(_11015_),
    .Y(_11032_));
 sky130_fd_sc_hd__a31o_2 _17735_ (.A1(_10986_),
    .A2(_10987_),
    .A3(_10988_),
    .B1(_10991_),
    .X(_11033_));
 sky130_fd_sc_hd__xor2_1 _17736_ (.A(_11011_),
    .B(_11033_),
    .X(_11034_));
 sky130_fd_sc_hd__or2_2 _17737_ (.A(_10972_),
    .B(_10974_),
    .X(_11035_));
 sky130_fd_sc_hd__buf_2 _17738_ (.A(_10968_),
    .X(_11036_));
 sky130_fd_sc_hd__buf_2 _17739_ (.A(_11036_),
    .X(_11037_));
 sky130_fd_sc_hd__buf_2 _17740_ (.A(_10976_),
    .X(_11038_));
 sky130_fd_sc_hd__clkbuf_4 _17741_ (.A(_11038_),
    .X(_11039_));
 sky130_fd_sc_hd__nand4_1 _17742_ (.A(_10641_),
    .B(_10612_),
    .C(_11037_),
    .D(_11039_),
    .Y(_11040_));
 sky130_fd_sc_hd__buf_2 _17743_ (.A(_10631_),
    .X(_11041_));
 sky130_fd_sc_hd__buf_2 _17744_ (.A(_10969_),
    .X(_11042_));
 sky130_fd_sc_hd__buf_2 _17745_ (.A(_11038_),
    .X(_11043_));
 sky130_fd_sc_hd__buf_2 _17746_ (.A(_10599_),
    .X(_11044_));
 sky130_fd_sc_hd__a22o_1 _17747_ (.A1(_11041_),
    .A2(_11042_),
    .B1(_11043_),
    .B2(_11044_),
    .X(_11045_));
 sky130_fd_sc_hd__nand2_1 _17748_ (.A(_11040_),
    .B(_11045_),
    .Y(_11046_));
 sky130_fd_sc_hd__clkbuf_2 _17749_ (.A(\genblk1.pcpi_mul.rs1[8] ),
    .X(_11047_));
 sky130_fd_sc_hd__buf_2 _17750_ (.A(_11047_),
    .X(_11048_));
 sky130_fd_sc_hd__clkbuf_4 _17751_ (.A(_11048_),
    .X(_11049_));
 sky130_fd_sc_hd__clkbuf_4 _17752_ (.A(_11049_),
    .X(_11050_));
 sky130_fd_sc_hd__nand2_1 _17753_ (.A(_10645_),
    .B(_11050_),
    .Y(_11051_));
 sky130_fd_sc_hd__xor2_1 _17754_ (.A(_11046_),
    .B(_11051_),
    .X(_11052_));
 sky130_fd_sc_hd__buf_2 _17755_ (.A(_10695_),
    .X(_11053_));
 sky130_fd_sc_hd__clkbuf_2 _17756_ (.A(\genblk1.pcpi_mul.rs1[11] ),
    .X(_11054_));
 sky130_fd_sc_hd__buf_2 _17757_ (.A(_11054_),
    .X(_11055_));
 sky130_fd_sc_hd__clkbuf_4 _17758_ (.A(_11055_),
    .X(_11056_));
 sky130_fd_sc_hd__buf_2 _17759_ (.A(_10670_),
    .X(_11057_));
 sky130_fd_sc_hd__clkbuf_2 _17760_ (.A(_10707_),
    .X(_11058_));
 sky130_fd_sc_hd__buf_2 _17761_ (.A(_10909_),
    .X(_11059_));
 sky130_fd_sc_hd__nand4_2 _17762_ (.A(_11057_),
    .B(_11058_),
    .C(_10912_),
    .D(_11059_),
    .Y(_11060_));
 sky130_fd_sc_hd__clkbuf_2 _17763_ (.A(_10701_),
    .X(_11061_));
 sky130_fd_sc_hd__buf_2 _17764_ (.A(_10909_),
    .X(_11062_));
 sky130_fd_sc_hd__buf_2 _17765_ (.A(_10661_),
    .X(_11063_));
 sky130_fd_sc_hd__a22o_1 _17766_ (.A1(_11061_),
    .A2(_10757_),
    .B1(_11062_),
    .B2(_11063_),
    .X(_11064_));
 sky130_fd_sc_hd__nand4_2 _17767_ (.A(_11053_),
    .B(_11056_),
    .C(_11060_),
    .D(_11064_),
    .Y(_11065_));
 sky130_fd_sc_hd__buf_2 _17768_ (.A(\genblk1.pcpi_mul.rs1[11] ),
    .X(_11066_));
 sky130_fd_sc_hd__buf_2 _17769_ (.A(_11066_),
    .X(_11067_));
 sky130_fd_sc_hd__clkbuf_4 _17770_ (.A(_11067_),
    .X(_11068_));
 sky130_fd_sc_hd__a22o_1 _17771_ (.A1(_10584_),
    .A2(_11068_),
    .B1(_11060_),
    .B2(_11064_),
    .X(_11069_));
 sky130_fd_sc_hd__o21bai_2 _17772_ (.A1(_10977_),
    .A2(_10980_),
    .B1_N(_10979_),
    .Y(_11070_));
 sky130_fd_sc_hd__nand3_1 _17773_ (.A(_11065_),
    .B(_11069_),
    .C(_11070_),
    .Y(_11071_));
 sky130_fd_sc_hd__a21o_1 _17774_ (.A1(_11065_),
    .A2(_11069_),
    .B1(_11070_),
    .X(_11072_));
 sky130_fd_sc_hd__nand3_1 _17775_ (.A(_11052_),
    .B(_11071_),
    .C(_11072_),
    .Y(_11073_));
 sky130_fd_sc_hd__a21o_1 _17776_ (.A1(_11071_),
    .A2(_11072_),
    .B1(_11052_),
    .X(_11074_));
 sky130_fd_sc_hd__a21bo_1 _17777_ (.A1(_10975_),
    .A2(_10985_),
    .B1_N(_10984_),
    .X(_11075_));
 sky130_fd_sc_hd__and3_2 _17778_ (.A(_11073_),
    .B(_11074_),
    .C(_11075_),
    .X(_11076_));
 sky130_fd_sc_hd__a21oi_2 _17779_ (.A1(_11073_),
    .A2(_11074_),
    .B1(_11075_),
    .Y(_11077_));
 sky130_fd_sc_hd__a211oi_4 _17780_ (.A1(_10970_),
    .A2(_11035_),
    .B1(_11076_),
    .C1(_11077_),
    .Y(_11078_));
 sky130_fd_sc_hd__o211a_1 _17781_ (.A1(_11076_),
    .A2(_11077_),
    .B1(_10970_),
    .C1(_11035_),
    .X(_11079_));
 sky130_fd_sc_hd__clkbuf_4 _17782_ (.A(_10737_),
    .X(_11080_));
 sky130_fd_sc_hd__a31o_1 _17783_ (.A1(_10667_),
    .A2(_11080_),
    .A3(_11000_),
    .B1(_10996_),
    .X(_11081_));
 sky130_fd_sc_hd__buf_2 _17784_ (.A(_10995_),
    .X(_11082_));
 sky130_fd_sc_hd__and4_1 _17785_ (.A(_10675_),
    .B(_10665_),
    .C(_11082_),
    .D(_10998_),
    .X(_11083_));
 sky130_fd_sc_hd__clkbuf_4 _17786_ (.A(_10995_),
    .X(_11084_));
 sky130_fd_sc_hd__buf_2 _17787_ (.A(\genblk1.pcpi_mul.rs2[8] ),
    .X(_11085_));
 sky130_fd_sc_hd__clkbuf_4 _17788_ (.A(_11085_),
    .X(_11086_));
 sky130_fd_sc_hd__clkbuf_2 _17789_ (.A(_10861_),
    .X(_11087_));
 sky130_fd_sc_hd__a22oi_1 _17790_ (.A1(_10742_),
    .A2(_11084_),
    .B1(_11086_),
    .B2(_11087_),
    .Y(_11088_));
 sky130_fd_sc_hd__clkbuf_2 _17791_ (.A(_10993_),
    .X(_11089_));
 sky130_fd_sc_hd__and4bb_1 _17792_ (.A_N(_11083_),
    .B_N(_11088_),
    .C(_11089_),
    .D(_10855_),
    .X(_11090_));
 sky130_fd_sc_hd__buf_2 _17793_ (.A(_10697_),
    .X(_11091_));
 sky130_fd_sc_hd__o2bb2a_1 _17794_ (.A1_N(_11089_),
    .A2_N(_11091_),
    .B1(_11083_),
    .B2(_11088_),
    .X(_11092_));
 sky130_fd_sc_hd__or3b_1 _17795_ (.A(_11090_),
    .B(_11092_),
    .C_N(_10965_),
    .X(_11093_));
 sky130_fd_sc_hd__o21bai_2 _17796_ (.A1(_11090_),
    .A2(_11092_),
    .B1_N(_10965_),
    .Y(_11094_));
 sky130_fd_sc_hd__and3_1 _17797_ (.A(_11081_),
    .B(_11093_),
    .C(_11094_),
    .X(_11095_));
 sky130_fd_sc_hd__a21oi_1 _17798_ (.A1(_11093_),
    .A2(_11094_),
    .B1(_11081_),
    .Y(_11096_));
 sky130_fd_sc_hd__or2_1 _17799_ (.A(_11095_),
    .B(_11096_),
    .X(_11097_));
 sky130_fd_sc_hd__nand2_1 _17800_ (.A(_11001_),
    .B(_11002_),
    .Y(_11098_));
 sky130_fd_sc_hd__o21a_1 _17801_ (.A1(_10901_),
    .A2(_11003_),
    .B1(_11098_),
    .X(_11099_));
 sky130_fd_sc_hd__xnor2_1 _17802_ (.A(_11097_),
    .B(_11099_),
    .Y(_11100_));
 sky130_fd_sc_hd__nor3_2 _17803_ (.A(_11078_),
    .B(_11079_),
    .C(_11100_),
    .Y(_11101_));
 sky130_fd_sc_hd__o21a_1 _17804_ (.A1(_11078_),
    .A2(_11079_),
    .B1(_11100_),
    .X(_11102_));
 sky130_fd_sc_hd__a211oi_4 _17805_ (.A1(_11007_),
    .A2(_11009_),
    .B1(_11101_),
    .C1(_11102_),
    .Y(_11103_));
 sky130_fd_sc_hd__o211a_1 _17806_ (.A1(_11101_),
    .A2(_11102_),
    .B1(_11007_),
    .C1(_11009_),
    .X(_11104_));
 sky130_fd_sc_hd__nand2_1 _17807_ (.A(_10609_),
    .B(_10895_),
    .Y(_11105_));
 sky130_fd_sc_hd__clkbuf_2 _17808_ (.A(\genblk1.pcpi_mul.rs2[11] ),
    .X(_11106_));
 sky130_fd_sc_hd__clkbuf_2 _17809_ (.A(_11106_),
    .X(_11107_));
 sky130_fd_sc_hd__clkbuf_4 _17810_ (.A(_11107_),
    .X(_11108_));
 sky130_fd_sc_hd__buf_4 _17811_ (.A(_11108_),
    .X(_11109_));
 sky130_fd_sc_hd__clkbuf_2 _17812_ (.A(\genblk1.pcpi_mul.rs2[11] ),
    .X(_11110_));
 sky130_fd_sc_hd__buf_2 _17813_ (.A(_11110_),
    .X(_11111_));
 sky130_fd_sc_hd__buf_2 _17814_ (.A(_11111_),
    .X(_11112_));
 sky130_fd_sc_hd__buf_2 _17815_ (.A(_10710_),
    .X(_11113_));
 sky130_fd_sc_hd__a22o_1 _17816_ (.A1(_10638_),
    .A2(_10957_),
    .B1(_11112_),
    .B2(_11113_),
    .X(_11114_));
 sky130_fd_sc_hd__a21bo_1 _17817_ (.A1(_11109_),
    .A2(_10964_),
    .B1_N(_11114_),
    .X(_11115_));
 sky130_fd_sc_hd__xor2_1 _17818_ (.A(_11105_),
    .B(_11115_),
    .X(_11116_));
 sky130_fd_sc_hd__nor3b_1 _17819_ (.A(_11103_),
    .B(_11104_),
    .C_N(_11116_),
    .Y(_11117_));
 sky130_fd_sc_hd__o21ba_1 _17820_ (.A1(_11103_),
    .A2(_11104_),
    .B1_N(_11116_),
    .X(_11118_));
 sky130_fd_sc_hd__or3_1 _17821_ (.A(_11013_),
    .B(net354),
    .C(_11118_),
    .X(_11119_));
 sky130_fd_sc_hd__o21ai_1 _17822_ (.A1(net354),
    .A2(_11118_),
    .B1(_11013_),
    .Y(_11120_));
 sky130_fd_sc_hd__nand3_1 _17823_ (.A(_11034_),
    .B(_11119_),
    .C(_11120_),
    .Y(_11121_));
 sky130_fd_sc_hd__a21o_1 _17824_ (.A1(_11119_),
    .A2(_11120_),
    .B1(_11034_),
    .X(_11122_));
 sky130_fd_sc_hd__o211a_1 _17825_ (.A1(_11032_),
    .A2(_11019_),
    .B1(_11121_),
    .C1(_11122_),
    .X(_11123_));
 sky130_fd_sc_hd__a211oi_1 _17826_ (.A1(_11121_),
    .A2(_11122_),
    .B1(_11032_),
    .C1(_11019_),
    .Y(_11124_));
 sky130_fd_sc_hd__nor3_1 _17827_ (.A(_11031_),
    .B(_11123_),
    .C(_11124_),
    .Y(_11125_));
 sky130_fd_sc_hd__o21a_1 _17828_ (.A1(_11123_),
    .A2(_11124_),
    .B1(_11031_),
    .X(_11126_));
 sky130_fd_sc_hd__a211oi_1 _17829_ (.A1(_11022_),
    .A2(_11025_),
    .B1(_11125_),
    .C1(_11126_),
    .Y(_11127_));
 sky130_fd_sc_hd__o211a_1 _17830_ (.A1(_11125_),
    .A2(_11126_),
    .B1(_11022_),
    .C1(_11025_),
    .X(_11128_));
 sky130_fd_sc_hd__or2_1 _17831_ (.A(_11127_),
    .B(_11128_),
    .X(_11129_));
 sky130_fd_sc_hd__nand3_1 _17832_ (.A(_11024_),
    .B(_11025_),
    .C(_11026_),
    .Y(_11130_));
 sky130_fd_sc_hd__a211o_1 _17833_ (.A1(_10954_),
    .A2(_10951_),
    .B1(_11027_),
    .C1(_11028_),
    .X(_11131_));
 sky130_fd_sc_hd__nand2_1 _17834_ (.A(_11130_),
    .B(_11131_),
    .Y(_11132_));
 sky130_fd_sc_hd__xnor2_1 _17835_ (.A(_11129_),
    .B(_11132_),
    .Y(_00057_));
 sky130_fd_sc_hd__nand2_1 _17836_ (.A(_11011_),
    .B(_11033_),
    .Y(_11133_));
 sky130_fd_sc_hd__clkbuf_2 _17837_ (.A(\genblk1.pcpi_mul.rs2[12] ),
    .X(_11134_));
 sky130_fd_sc_hd__clkbuf_4 _17838_ (.A(_11134_),
    .X(_11135_));
 sky130_fd_sc_hd__clkbuf_2 _17839_ (.A(_11135_),
    .X(_11136_));
 sky130_fd_sc_hd__buf_4 _17840_ (.A(_11136_),
    .X(_11137_));
 sky130_fd_sc_hd__clkbuf_4 _17841_ (.A(_10961_),
    .X(_11138_));
 sky130_fd_sc_hd__nand2_1 _17842_ (.A(_10651_),
    .B(_11138_),
    .Y(_11139_));
 sky130_fd_sc_hd__clkbuf_2 _17843_ (.A(\genblk1.pcpi_mul.rs2[10] ),
    .X(_11140_));
 sky130_fd_sc_hd__clkbuf_2 _17844_ (.A(_11140_),
    .X(_11141_));
 sky130_fd_sc_hd__buf_2 _17845_ (.A(_11141_),
    .X(_11142_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17846_ (.A(\genblk1.pcpi_mul.rs2[11] ),
    .X(_11143_));
 sky130_fd_sc_hd__clkbuf_2 _17847_ (.A(_11143_),
    .X(_11144_));
 sky130_fd_sc_hd__buf_2 _17848_ (.A(_11144_),
    .X(_11145_));
 sky130_fd_sc_hd__and4_1 _17849_ (.A(_10595_),
    .B(_10629_),
    .C(_11142_),
    .D(_11145_),
    .X(_11146_));
 sky130_fd_sc_hd__a22o_1 _17850_ (.A1(_10629_),
    .A2(_11142_),
    .B1(_11108_),
    .B2(_10595_),
    .X(_11147_));
 sky130_fd_sc_hd__and2b_1 _17851_ (.A_N(_11146_),
    .B(_11147_),
    .X(_11148_));
 sky130_fd_sc_hd__xnor2_1 _17852_ (.A(_11139_),
    .B(_11148_),
    .Y(_11149_));
 sky130_fd_sc_hd__and3_1 _17853_ (.A(_10590_),
    .B(_11137_),
    .C(_11149_),
    .X(_11150_));
 sky130_fd_sc_hd__a21oi_1 _17854_ (.A1(_10603_),
    .A2(_11137_),
    .B1(_11149_),
    .Y(_11151_));
 sky130_fd_sc_hd__nor2_1 _17855_ (.A(_11150_),
    .B(_11151_),
    .Y(_11152_));
 sky130_fd_sc_hd__o21a_1 _17856_ (.A1(_11046_),
    .A2(_11051_),
    .B1(_11040_),
    .X(_11153_));
 sky130_fd_sc_hd__buf_2 _17857_ (.A(\genblk1.pcpi_mul.rs1[10] ),
    .X(_11154_));
 sky130_fd_sc_hd__buf_2 _17858_ (.A(_11154_),
    .X(_11155_));
 sky130_fd_sc_hd__buf_2 _17859_ (.A(_11155_),
    .X(_11156_));
 sky130_fd_sc_hd__buf_4 _17860_ (.A(_11156_),
    .X(_11157_));
 sky130_fd_sc_hd__nand2_1 _17861_ (.A(_10612_),
    .B(_11157_),
    .Y(_11158_));
 sky130_fd_sc_hd__buf_2 _17862_ (.A(\genblk1.pcpi_mul.rs1[11] ),
    .X(_11159_));
 sky130_fd_sc_hd__buf_2 _17863_ (.A(_11159_),
    .X(_11160_));
 sky130_fd_sc_hd__buf_4 _17864_ (.A(_11160_),
    .X(_11161_));
 sky130_fd_sc_hd__nand2_1 _17865_ (.A(_10627_),
    .B(_11161_),
    .Y(_11162_));
 sky130_fd_sc_hd__nand2_1 _17866_ (.A(_10641_),
    .B(_11039_),
    .Y(_11163_));
 sky130_fd_sc_hd__nand2_1 _17867_ (.A(_10632_),
    .B(_11056_),
    .Y(_11164_));
 sky130_fd_sc_hd__nor2_1 _17868_ (.A(_11163_),
    .B(_11164_),
    .Y(_11165_));
 sky130_fd_sc_hd__a21oi_1 _17869_ (.A1(_11158_),
    .A2(_11162_),
    .B1(_11165_),
    .Y(_11166_));
 sky130_fd_sc_hd__buf_4 _17870_ (.A(_11042_),
    .X(_11167_));
 sky130_fd_sc_hd__nand2_1 _17871_ (.A(_10645_),
    .B(_11167_),
    .Y(_11168_));
 sky130_fd_sc_hd__xnor2_1 _17872_ (.A(_11166_),
    .B(_11168_),
    .Y(_11169_));
 sky130_fd_sc_hd__buf_2 _17873_ (.A(\genblk1.pcpi_mul.rs1[12] ),
    .X(_11170_));
 sky130_fd_sc_hd__clkbuf_2 _17874_ (.A(_11170_),
    .X(_11171_));
 sky130_fd_sc_hd__clkbuf_4 _17875_ (.A(_11171_),
    .X(_11172_));
 sky130_fd_sc_hd__nand2_1 _17876_ (.A(_11053_),
    .B(_11172_),
    .Y(_11173_));
 sky130_fd_sc_hd__buf_2 _17877_ (.A(\genblk1.pcpi_mul.rs1[8] ),
    .X(_11174_));
 sky130_fd_sc_hd__clkbuf_2 _17878_ (.A(_11174_),
    .X(_11175_));
 sky130_fd_sc_hd__and4_1 _17879_ (.A(_11063_),
    .B(_10708_),
    .C(_11062_),
    .D(_11175_),
    .X(_11176_));
 sky130_fd_sc_hd__clkbuf_4 _17880_ (.A(_10967_),
    .X(_11177_));
 sky130_fd_sc_hd__a22oi_2 _17881_ (.A1(_11058_),
    .A2(_11059_),
    .B1(_11177_),
    .B2(_10662_),
    .Y(_11178_));
 sky130_fd_sc_hd__nor2_1 _17882_ (.A(_11176_),
    .B(_11178_),
    .Y(_11179_));
 sky130_fd_sc_hd__xnor2_1 _17883_ (.A(_11173_),
    .B(_11179_),
    .Y(_11180_));
 sky130_fd_sc_hd__and2_1 _17884_ (.A(_11060_),
    .B(_11065_),
    .X(_11181_));
 sky130_fd_sc_hd__xnor2_1 _17885_ (.A(_11180_),
    .B(_11181_),
    .Y(_11182_));
 sky130_fd_sc_hd__xnor2_1 _17886_ (.A(_11169_),
    .B(_11182_),
    .Y(_11183_));
 sky130_fd_sc_hd__and2_1 _17887_ (.A(_11071_),
    .B(_11073_),
    .X(_11184_));
 sky130_fd_sc_hd__xor2_1 _17888_ (.A(_11183_),
    .B(_11184_),
    .X(_11185_));
 sky130_fd_sc_hd__xnor2_1 _17889_ (.A(_11153_),
    .B(_11185_),
    .Y(_11186_));
 sky130_fd_sc_hd__nor2_1 _17890_ (.A(_11098_),
    .B(_11097_),
    .Y(_11187_));
 sky130_fd_sc_hd__or2_1 _17891_ (.A(_11083_),
    .B(_11090_),
    .X(_11188_));
 sky130_fd_sc_hd__clkbuf_2 _17892_ (.A(\genblk1.pcpi_mul.rs2[9] ),
    .X(_11189_));
 sky130_fd_sc_hd__clkbuf_2 _17893_ (.A(_11189_),
    .X(_11190_));
 sky130_fd_sc_hd__clkbuf_4 _17894_ (.A(_11190_),
    .X(_11191_));
 sky130_fd_sc_hd__a32o_1 _17895_ (.A1(_10630_),
    .A2(_11191_),
    .A3(_11114_),
    .B1(_10964_),
    .B2(_11109_),
    .X(_11192_));
 sky130_fd_sc_hd__buf_2 _17896_ (.A(_10757_),
    .X(_11193_));
 sky130_fd_sc_hd__nand2_1 _17897_ (.A(_10737_),
    .B(_11193_),
    .Y(_11194_));
 sky130_fd_sc_hd__buf_2 _17898_ (.A(\genblk1.pcpi_mul.rs2[8] ),
    .X(_11195_));
 sky130_fd_sc_hd__clkbuf_2 _17899_ (.A(_11195_),
    .X(_11196_));
 sky130_fd_sc_hd__clkbuf_4 _17900_ (.A(_11196_),
    .X(_11197_));
 sky130_fd_sc_hd__nand4_2 _17901_ (.A(_10797_),
    .B(_10855_),
    .C(_10783_),
    .D(_11197_),
    .Y(_11198_));
 sky130_fd_sc_hd__buf_2 _17902_ (.A(_10790_),
    .X(_11199_));
 sky130_fd_sc_hd__clkbuf_2 _17903_ (.A(_10839_),
    .X(_11200_));
 sky130_fd_sc_hd__clkbuf_4 _17904_ (.A(_11200_),
    .X(_11201_));
 sky130_fd_sc_hd__a22o_1 _17905_ (.A1(_11199_),
    .A2(_11084_),
    .B1(_11201_),
    .B2(_10797_),
    .X(_11202_));
 sky130_fd_sc_hd__nand3b_1 _17906_ (.A_N(_11194_),
    .B(_11198_),
    .C(_11202_),
    .Y(_11203_));
 sky130_fd_sc_hd__a21bo_1 _17907_ (.A1(_11198_),
    .A2(_11202_),
    .B1_N(_11194_),
    .X(_11204_));
 sky130_fd_sc_hd__nand2_1 _17908_ (.A(_11203_),
    .B(_11204_),
    .Y(_11205_));
 sky130_fd_sc_hd__xnor2_1 _17909_ (.A(_11192_),
    .B(_11205_),
    .Y(_11206_));
 sky130_fd_sc_hd__xor2_1 _17910_ (.A(_11188_),
    .B(_11206_),
    .X(_11207_));
 sky130_fd_sc_hd__a21boi_2 _17911_ (.A1(_11081_),
    .A2(_11094_),
    .B1_N(_11093_),
    .Y(_11208_));
 sky130_fd_sc_hd__xnor2_1 _17912_ (.A(_11207_),
    .B(_11208_),
    .Y(_11209_));
 sky130_fd_sc_hd__xor2_1 _17913_ (.A(_11187_),
    .B(_11209_),
    .X(_11210_));
 sky130_fd_sc_hd__xnor2_1 _17914_ (.A(_11186_),
    .B(_11210_),
    .Y(_11211_));
 sky130_fd_sc_hd__nor2_1 _17915_ (.A(_11003_),
    .B(_11097_),
    .Y(_11212_));
 sky130_fd_sc_hd__a21o_1 _17916_ (.A1(_11004_),
    .A2(_11212_),
    .B1(_11101_),
    .X(_11213_));
 sky130_fd_sc_hd__xnor2_1 _17917_ (.A(_11211_),
    .B(_11213_),
    .Y(_11214_));
 sky130_fd_sc_hd__xnor2_1 _17918_ (.A(_11152_),
    .B(_11214_),
    .Y(_11215_));
 sky130_fd_sc_hd__xnor2_1 _17919_ (.A(_11117_),
    .B(_11215_),
    .Y(_11216_));
 sky130_fd_sc_hd__o21ai_1 _17920_ (.A1(_11076_),
    .A2(_11078_),
    .B1(_11103_),
    .Y(_11217_));
 sky130_fd_sc_hd__or3_1 _17921_ (.A(_11076_),
    .B(_11078_),
    .C(_11103_),
    .X(_11218_));
 sky130_fd_sc_hd__and2_1 _17922_ (.A(_11217_),
    .B(_11218_),
    .X(_11219_));
 sky130_fd_sc_hd__xnor2_1 _17923_ (.A(_11216_),
    .B(_11219_),
    .Y(_11220_));
 sky130_fd_sc_hd__nand2_1 _17924_ (.A(_11119_),
    .B(_11121_),
    .Y(_11221_));
 sky130_fd_sc_hd__xnor2_1 _17925_ (.A(_11220_),
    .B(_11221_),
    .Y(_11222_));
 sky130_fd_sc_hd__xor2_1 _17926_ (.A(_11133_),
    .B(_11222_),
    .X(_11223_));
 sky130_fd_sc_hd__nor2_1 _17927_ (.A(_11123_),
    .B(_11125_),
    .Y(_11224_));
 sky130_fd_sc_hd__xnor2_1 _17928_ (.A(_11223_),
    .B(_11224_),
    .Y(_11225_));
 sky130_vsdinv _17929_ (.A(_11127_),
    .Y(_11226_));
 sky130_fd_sc_hd__a31oi_1 _17930_ (.A1(_11130_),
    .A2(_11131_),
    .A3(_11226_),
    .B1(_11128_),
    .Y(_11227_));
 sky130_fd_sc_hd__xnor2_1 _17931_ (.A(_11225_),
    .B(_11227_),
    .Y(_00058_));
 sky130_fd_sc_hd__or2b_1 _17932_ (.A(_11220_),
    .B_N(_11221_),
    .X(_11228_));
 sky130_fd_sc_hd__or2b_1 _17933_ (.A(_11133_),
    .B_N(_11222_),
    .X(_11229_));
 sky130_fd_sc_hd__or4b_1 _17934_ (.A(_11103_),
    .B(_11104_),
    .C(_11215_),
    .D_N(_11116_),
    .X(_11230_));
 sky130_fd_sc_hd__nand2_1 _17935_ (.A(_11216_),
    .B(_11219_),
    .Y(_11231_));
 sky130_fd_sc_hd__and2_1 _17936_ (.A(_11152_),
    .B(_11214_),
    .X(_11232_));
 sky130_fd_sc_hd__buf_2 _17937_ (.A(_11135_),
    .X(_11233_));
 sky130_fd_sc_hd__buf_2 _17938_ (.A(\genblk1.pcpi_mul.rs2[13] ),
    .X(_11234_));
 sky130_fd_sc_hd__buf_2 _17939_ (.A(_11234_),
    .X(_11235_));
 sky130_fd_sc_hd__buf_2 _17940_ (.A(_11235_),
    .X(_11236_));
 sky130_fd_sc_hd__buf_4 _17941_ (.A(_11236_),
    .X(_11237_));
 sky130_fd_sc_hd__a22oi_1 _17942_ (.A1(_10596_),
    .A2(_11233_),
    .B1(_11237_),
    .B2(_10623_),
    .Y(_11238_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17943_ (.A(\genblk1.pcpi_mul.rs2[13] ),
    .X(_11239_));
 sky130_fd_sc_hd__buf_1 _17944_ (.A(_11239_),
    .X(_11240_));
 sky130_fd_sc_hd__clkbuf_4 _17945_ (.A(_11240_),
    .X(_11241_));
 sky130_fd_sc_hd__buf_2 _17946_ (.A(_11241_),
    .X(_11242_));
 sky130_fd_sc_hd__and4_1 _17947_ (.A(_10589_),
    .B(_10636_),
    .C(_11135_),
    .D(_11242_),
    .X(_11243_));
 sky130_fd_sc_hd__nor2_1 _17948_ (.A(_11238_),
    .B(_11243_),
    .Y(_11244_));
 sky130_fd_sc_hd__buf_2 _17949_ (.A(_10797_),
    .X(_11245_));
 sky130_fd_sc_hd__nand2_1 _17950_ (.A(_11245_),
    .B(_11138_),
    .Y(_11246_));
 sky130_fd_sc_hd__and4_1 _17951_ (.A(_10629_),
    .B(_11087_),
    .C(_10957_),
    .D(_11145_),
    .X(_11247_));
 sky130_fd_sc_hd__a22o_1 _17952_ (.A1(_11087_),
    .A2(_10957_),
    .B1(_11108_),
    .B2(_10629_),
    .X(_11248_));
 sky130_fd_sc_hd__and2b_1 _17953_ (.A_N(_11247_),
    .B(_11248_),
    .X(_11249_));
 sky130_fd_sc_hd__xnor2_1 _17954_ (.A(_11246_),
    .B(_11249_),
    .Y(_11250_));
 sky130_fd_sc_hd__and2_1 _17955_ (.A(_11244_),
    .B(_11250_),
    .X(_11251_));
 sky130_fd_sc_hd__nor2_1 _17956_ (.A(_11244_),
    .B(_11250_),
    .Y(_11252_));
 sky130_fd_sc_hd__or2_1 _17957_ (.A(_11251_),
    .B(_11252_),
    .X(_11253_));
 sky130_fd_sc_hd__nand2_1 _17958_ (.A(_11187_),
    .B(_11209_),
    .Y(_11254_));
 sky130_fd_sc_hd__nand2_1 _17959_ (.A(_11186_),
    .B(_11210_),
    .Y(_11255_));
 sky130_fd_sc_hd__or2_1 _17960_ (.A(_11163_),
    .B(_11164_),
    .X(_11256_));
 sky130_fd_sc_hd__a211o_1 _17961_ (.A1(_11158_),
    .A2(_11162_),
    .B1(_11165_),
    .C1(_11168_),
    .X(_11257_));
 sky130_fd_sc_hd__or2b_1 _17962_ (.A(_11181_),
    .B_N(_11180_),
    .X(_11258_));
 sky130_fd_sc_hd__nand2_1 _17963_ (.A(_11169_),
    .B(_11182_),
    .Y(_11259_));
 sky130_fd_sc_hd__buf_2 _17964_ (.A(\genblk1.pcpi_mul.rs1[12] ),
    .X(_11260_));
 sky130_fd_sc_hd__buf_2 _17965_ (.A(_11260_),
    .X(_11261_));
 sky130_fd_sc_hd__clkbuf_4 _17966_ (.A(_11261_),
    .X(_11262_));
 sky130_fd_sc_hd__nand2_1 _17967_ (.A(_10627_),
    .B(_11262_),
    .Y(_11263_));
 sky130_fd_sc_hd__clkbuf_4 _17968_ (.A(_11067_),
    .X(_11264_));
 sky130_fd_sc_hd__clkbuf_4 _17969_ (.A(_11171_),
    .X(_11265_));
 sky130_fd_sc_hd__and4_1 _17970_ (.A(_11044_),
    .B(_11041_),
    .C(_11264_),
    .D(_11265_),
    .X(_11266_));
 sky130_fd_sc_hd__a21oi_1 _17971_ (.A1(_11164_),
    .A2(_11263_),
    .B1(_11266_),
    .Y(_11267_));
 sky130_fd_sc_hd__buf_2 _17972_ (.A(\genblk1.pcpi_mul.rs1[10] ),
    .X(_11268_));
 sky130_fd_sc_hd__clkbuf_4 _17973_ (.A(_11268_),
    .X(_11269_));
 sky130_fd_sc_hd__buf_2 _17974_ (.A(_11269_),
    .X(_11270_));
 sky130_fd_sc_hd__and2_1 _17975_ (.A(_10625_),
    .B(_11270_),
    .X(_11271_));
 sky130_fd_sc_hd__nor2_1 _17976_ (.A(_11267_),
    .B(_11271_),
    .Y(_11272_));
 sky130_fd_sc_hd__and2_1 _17977_ (.A(_11267_),
    .B(_11271_),
    .X(_11273_));
 sky130_fd_sc_hd__nor2_1 _17978_ (.A(_11272_),
    .B(_11273_),
    .Y(_11274_));
 sky130_fd_sc_hd__clkbuf_2 _17979_ (.A(\genblk1.pcpi_mul.rs1[13] ),
    .X(_11275_));
 sky130_fd_sc_hd__clkbuf_4 _17980_ (.A(_11275_),
    .X(_11276_));
 sky130_fd_sc_hd__clkbuf_4 _17981_ (.A(_11276_),
    .X(_11277_));
 sky130_fd_sc_hd__buf_2 _17982_ (.A(_11277_),
    .X(_11278_));
 sky130_fd_sc_hd__nand2_1 _17983_ (.A(_10584_),
    .B(_11278_),
    .Y(_11279_));
 sky130_fd_sc_hd__buf_2 _17984_ (.A(_10968_),
    .X(_11280_));
 sky130_fd_sc_hd__and4_1 _17985_ (.A(_11057_),
    .B(_11058_),
    .C(_11175_),
    .D(_11280_),
    .X(_11281_));
 sky130_fd_sc_hd__buf_2 _17986_ (.A(_10708_),
    .X(_11282_));
 sky130_fd_sc_hd__a22oi_1 _17987_ (.A1(_11282_),
    .A2(_11049_),
    .B1(_11042_),
    .B2(_10662_),
    .Y(_11283_));
 sky130_fd_sc_hd__nor2_1 _17988_ (.A(_11281_),
    .B(_11283_),
    .Y(_11284_));
 sky130_fd_sc_hd__xnor2_2 _17989_ (.A(_11279_),
    .B(_11284_),
    .Y(_11285_));
 sky130_fd_sc_hd__o21ba_1 _17990_ (.A1(_11173_),
    .A2(_11178_),
    .B1_N(_11176_),
    .X(_11286_));
 sky130_fd_sc_hd__xnor2_1 _17991_ (.A(_11285_),
    .B(_11286_),
    .Y(_11287_));
 sky130_fd_sc_hd__xnor2_1 _17992_ (.A(_11274_),
    .B(_11287_),
    .Y(_11288_));
 sky130_fd_sc_hd__a21oi_1 _17993_ (.A1(_11258_),
    .A2(_11259_),
    .B1(_11288_),
    .Y(_11289_));
 sky130_fd_sc_hd__and3_1 _17994_ (.A(_11258_),
    .B(_11259_),
    .C(_11288_),
    .X(_11290_));
 sky130_fd_sc_hd__a211oi_2 _17995_ (.A1(_11256_),
    .A2(_11257_),
    .B1(_11289_),
    .C1(_11290_),
    .Y(_11291_));
 sky130_fd_sc_hd__o211a_1 _17996_ (.A1(_11289_),
    .A2(_11290_),
    .B1(_11256_),
    .C1(_11257_),
    .X(_11292_));
 sky130_fd_sc_hd__or2b_1 _17997_ (.A(_11208_),
    .B_N(_11207_),
    .X(_11293_));
 sky130_fd_sc_hd__a32o_1 _17998_ (.A1(_11192_),
    .A2(_11203_),
    .A3(_11204_),
    .B1(_11206_),
    .B2(_11188_),
    .X(_11294_));
 sky130_fd_sc_hd__nand2_1 _17999_ (.A(_11198_),
    .B(_11203_),
    .Y(_11295_));
 sky130_fd_sc_hd__a31o_1 _18000_ (.A1(_10676_),
    .A2(_11191_),
    .A3(_11147_),
    .B1(_11146_),
    .X(_11296_));
 sky130_fd_sc_hd__clkbuf_4 _18001_ (.A(_10973_),
    .X(_11297_));
 sky130_fd_sc_hd__buf_2 _18002_ (.A(_10836_),
    .X(_11298_));
 sky130_fd_sc_hd__clkbuf_4 _18003_ (.A(_11298_),
    .X(_11299_));
 sky130_fd_sc_hd__nand4_2 _18004_ (.A(_11193_),
    .B(_11091_),
    .C(_11299_),
    .D(_11197_),
    .Y(_11300_));
 sky130_fd_sc_hd__clkbuf_2 _18005_ (.A(_10978_),
    .X(_11301_));
 sky130_fd_sc_hd__buf_2 _18006_ (.A(_11301_),
    .X(_11302_));
 sky130_fd_sc_hd__a22o_1 _18007_ (.A1(_11302_),
    .A2(_10783_),
    .B1(_11201_),
    .B2(_10855_),
    .X(_11303_));
 sky130_fd_sc_hd__nand4_2 _18008_ (.A(_11080_),
    .B(_11297_),
    .C(_11300_),
    .D(_11303_),
    .Y(_11304_));
 sky130_fd_sc_hd__a22o_1 _18009_ (.A1(_10737_),
    .A2(_11297_),
    .B1(_11300_),
    .B2(_11303_),
    .X(_11305_));
 sky130_fd_sc_hd__nand3_2 _18010_ (.A(_11296_),
    .B(_11304_),
    .C(_11305_),
    .Y(_11306_));
 sky130_fd_sc_hd__a21o_1 _18011_ (.A1(_11304_),
    .A2(_11305_),
    .B1(_11296_),
    .X(_11307_));
 sky130_fd_sc_hd__nand3_2 _18012_ (.A(_11295_),
    .B(_11306_),
    .C(_11307_),
    .Y(_11308_));
 sky130_fd_sc_hd__a21o_1 _18013_ (.A1(_11306_),
    .A2(_11307_),
    .B1(_11295_),
    .X(_11309_));
 sky130_fd_sc_hd__nand3_2 _18014_ (.A(_11150_),
    .B(_11308_),
    .C(_11309_),
    .Y(_11310_));
 sky130_fd_sc_hd__a21o_1 _18015_ (.A1(_11308_),
    .A2(_11309_),
    .B1(_11150_),
    .X(_11311_));
 sky130_fd_sc_hd__and3_1 _18016_ (.A(_11294_),
    .B(_11310_),
    .C(_11311_),
    .X(_11312_));
 sky130_fd_sc_hd__a21oi_1 _18017_ (.A1(_11310_),
    .A2(_11311_),
    .B1(_11294_),
    .Y(_11313_));
 sky130_fd_sc_hd__nor3_1 _18018_ (.A(_11293_),
    .B(_11312_),
    .C(_11313_),
    .Y(_11314_));
 sky130_fd_sc_hd__o21a_1 _18019_ (.A1(_11312_),
    .A2(_11313_),
    .B1(_11293_),
    .X(_11315_));
 sky130_fd_sc_hd__nor4_1 _18020_ (.A(_11291_),
    .B(_11292_),
    .C(_11314_),
    .D(_11315_),
    .Y(_11316_));
 sky130_fd_sc_hd__o22a_1 _18021_ (.A1(_11291_),
    .A2(_11292_),
    .B1(_11314_),
    .B2(_11315_),
    .X(_11317_));
 sky130_fd_sc_hd__a211oi_2 _18022_ (.A1(_11254_),
    .A2(_11255_),
    .B1(net353),
    .C1(_11317_),
    .Y(_11318_));
 sky130_fd_sc_hd__o211a_1 _18023_ (.A1(_11316_),
    .A2(_11317_),
    .B1(_11254_),
    .C1(_11255_),
    .X(_11319_));
 sky130_fd_sc_hd__or3_1 _18024_ (.A(_11253_),
    .B(_11318_),
    .C(_11319_),
    .X(_11320_));
 sky130_fd_sc_hd__o21ai_1 _18025_ (.A1(_11318_),
    .A2(_11319_),
    .B1(_11253_),
    .Y(_11321_));
 sky130_fd_sc_hd__and3_1 _18026_ (.A(_11232_),
    .B(_11320_),
    .C(_11321_),
    .X(_11322_));
 sky130_fd_sc_hd__a21oi_1 _18027_ (.A1(_11320_),
    .A2(_11321_),
    .B1(_11232_),
    .Y(_11323_));
 sky130_fd_sc_hd__and2b_1 _18028_ (.A_N(_11211_),
    .B(_11213_),
    .X(_11324_));
 sky130_fd_sc_hd__and2b_1 _18029_ (.A_N(_11153_),
    .B(_11185_),
    .X(_11325_));
 sky130_fd_sc_hd__o21bai_2 _18030_ (.A1(_11183_),
    .A2(_11184_),
    .B1_N(_11325_),
    .Y(_11326_));
 sky130_fd_sc_hd__xnor2_1 _18031_ (.A(_11324_),
    .B(_11326_),
    .Y(_11327_));
 sky130_fd_sc_hd__nor3_1 _18032_ (.A(_11322_),
    .B(_11323_),
    .C(_11327_),
    .Y(_11328_));
 sky130_fd_sc_hd__o21a_1 _18033_ (.A1(_11322_),
    .A2(_11323_),
    .B1(_11327_),
    .X(_11329_));
 sky130_fd_sc_hd__a211oi_1 _18034_ (.A1(_11230_),
    .A2(_11231_),
    .B1(_11328_),
    .C1(_11329_),
    .Y(_11330_));
 sky130_fd_sc_hd__o211a_1 _18035_ (.A1(_11328_),
    .A2(_11329_),
    .B1(_11230_),
    .C1(_11231_),
    .X(_11331_));
 sky130_fd_sc_hd__nor3_1 _18036_ (.A(_11217_),
    .B(_11330_),
    .C(_11331_),
    .Y(_11332_));
 sky130_fd_sc_hd__o21a_1 _18037_ (.A1(_11330_),
    .A2(_11331_),
    .B1(_11217_),
    .X(_11333_));
 sky130_fd_sc_hd__a211o_1 _18038_ (.A1(_11228_),
    .A2(_11229_),
    .B1(_11332_),
    .C1(_11333_),
    .X(_11334_));
 sky130_fd_sc_hd__o211ai_1 _18039_ (.A1(_11332_),
    .A2(_11333_),
    .B1(_11228_),
    .C1(_11229_),
    .Y(_11335_));
 sky130_fd_sc_hd__nand2_1 _18040_ (.A(_11334_),
    .B(_11335_),
    .Y(_11336_));
 sky130_fd_sc_hd__or2_1 _18041_ (.A(_11223_),
    .B(_11224_),
    .X(_11337_));
 sky130_fd_sc_hd__a311o_1 _18042_ (.A1(_11130_),
    .A2(_11131_),
    .A3(_11226_),
    .B1(_11128_),
    .C1(_11225_),
    .X(_11338_));
 sky130_fd_sc_hd__nand2_1 _18043_ (.A(_11337_),
    .B(_11338_),
    .Y(_11339_));
 sky130_fd_sc_hd__xnor2_1 _18044_ (.A(_11336_),
    .B(_11339_),
    .Y(_00059_));
 sky130_fd_sc_hd__and2_1 _18045_ (.A(_11324_),
    .B(_11326_),
    .X(_11340_));
 sky130_fd_sc_hd__nor2_1 _18046_ (.A(_11289_),
    .B(_11291_),
    .Y(_11341_));
 sky130_fd_sc_hd__xnor2_1 _18047_ (.A(_11318_),
    .B(_11341_),
    .Y(_11342_));
 sky130_fd_sc_hd__clkbuf_4 _18048_ (.A(_11199_),
    .X(_11343_));
 sky130_fd_sc_hd__nand2_1 _18049_ (.A(_11343_),
    .B(_11191_),
    .Y(_11344_));
 sky130_fd_sc_hd__and4_1 _18050_ (.A(_11087_),
    .B(_10721_),
    .C(_10963_),
    .D(_11111_),
    .X(_11345_));
 sky130_fd_sc_hd__a22o_1 _18051_ (.A1(_10721_),
    .A2(_11142_),
    .B1(_11145_),
    .B2(_11087_),
    .X(_11346_));
 sky130_fd_sc_hd__and2b_1 _18052_ (.A_N(_11345_),
    .B(_11346_),
    .X(_11347_));
 sky130_fd_sc_hd__xnor2_2 _18053_ (.A(_11344_),
    .B(_11347_),
    .Y(_11348_));
 sky130_fd_sc_hd__clkbuf_2 _18054_ (.A(\genblk1.pcpi_mul.rs2[12] ),
    .X(_11349_));
 sky130_fd_sc_hd__buf_2 _18055_ (.A(_11349_),
    .X(_11350_));
 sky130_fd_sc_hd__and2_1 _18056_ (.A(_10607_),
    .B(_11350_),
    .X(_11351_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18057_ (.A(\genblk1.pcpi_mul.rs2[14] ),
    .X(_11352_));
 sky130_fd_sc_hd__buf_4 _18058_ (.A(_11352_),
    .X(_11353_));
 sky130_fd_sc_hd__buf_4 _18059_ (.A(_11353_),
    .X(_11354_));
 sky130_fd_sc_hd__nand4_2 _18060_ (.A(_10710_),
    .B(_10705_),
    .C(_11241_),
    .D(_11354_),
    .Y(_11355_));
 sky130_fd_sc_hd__clkbuf_4 _18061_ (.A(_11234_),
    .X(_11356_));
 sky130_fd_sc_hd__a22o_1 _18062_ (.A1(_10786_),
    .A2(_11356_),
    .B1(_11354_),
    .B2(_10587_),
    .X(_11357_));
 sky130_fd_sc_hd__nand3_1 _18063_ (.A(_11351_),
    .B(_11355_),
    .C(_11357_),
    .Y(_11358_));
 sky130_fd_sc_hd__a21o_1 _18064_ (.A1(_11355_),
    .A2(_11357_),
    .B1(_11351_),
    .X(_11359_));
 sky130_fd_sc_hd__and3_1 _18065_ (.A(_11243_),
    .B(_11358_),
    .C(_11359_),
    .X(_11360_));
 sky130_fd_sc_hd__a21o_1 _18066_ (.A1(_11358_),
    .A2(_11359_),
    .B1(_11243_),
    .X(_11361_));
 sky130_fd_sc_hd__or2b_1 _18067_ (.A(_11360_),
    .B_N(_11361_),
    .X(_11362_));
 sky130_fd_sc_hd__xor2_2 _18068_ (.A(_11348_),
    .B(_11362_),
    .X(_11363_));
 sky130_vsdinv _18069_ (.A(_11314_),
    .Y(_11364_));
 sky130_fd_sc_hd__or4_1 _18070_ (.A(_11291_),
    .B(_11292_),
    .C(_11314_),
    .D(_11315_),
    .X(_11365_));
 sky130_fd_sc_hd__or2b_1 _18071_ (.A(_11286_),
    .B_N(_11285_),
    .X(_11366_));
 sky130_fd_sc_hd__nand2_1 _18072_ (.A(_11274_),
    .B(_11287_),
    .Y(_11367_));
 sky130_fd_sc_hd__clkbuf_4 _18073_ (.A(_10645_),
    .X(_11368_));
 sky130_fd_sc_hd__buf_4 _18074_ (.A(_11277_),
    .X(_11369_));
 sky130_fd_sc_hd__a22oi_1 _18075_ (.A1(_10633_),
    .A2(_11262_),
    .B1(_11369_),
    .B2(_10601_),
    .Y(_11370_));
 sky130_fd_sc_hd__clkbuf_2 _18076_ (.A(\genblk1.pcpi_mul.rs1[13] ),
    .X(_11371_));
 sky130_fd_sc_hd__buf_2 _18077_ (.A(_11371_),
    .X(_11372_));
 sky130_fd_sc_hd__buf_2 _18078_ (.A(_11372_),
    .X(_11373_));
 sky130_fd_sc_hd__and4_1 _18079_ (.A(_10627_),
    .B(_10612_),
    .C(_11172_),
    .D(_11373_),
    .X(_11374_));
 sky130_fd_sc_hd__nor2_1 _18080_ (.A(_11370_),
    .B(_11374_),
    .Y(_11375_));
 sky130_fd_sc_hd__a21oi_1 _18081_ (.A1(_11368_),
    .A2(_11161_),
    .B1(_11375_),
    .Y(_11376_));
 sky130_fd_sc_hd__and3_1 _18082_ (.A(_10680_),
    .B(_11161_),
    .C(_11375_),
    .X(_11377_));
 sky130_fd_sc_hd__nor2_1 _18083_ (.A(_11376_),
    .B(_11377_),
    .Y(_11378_));
 sky130_fd_sc_hd__buf_2 _18084_ (.A(\genblk1.pcpi_mul.rs1[14] ),
    .X(_11379_));
 sky130_fd_sc_hd__buf_2 _18085_ (.A(_11379_),
    .X(_11380_));
 sky130_fd_sc_hd__clkbuf_2 _18086_ (.A(_11380_),
    .X(_11381_));
 sky130_fd_sc_hd__buf_4 _18087_ (.A(_11381_),
    .X(_11382_));
 sky130_fd_sc_hd__nand2_1 _18088_ (.A(_10584_),
    .B(_11382_),
    .Y(_11383_));
 sky130_fd_sc_hd__and4_1 _18089_ (.A(_10672_),
    .B(_11282_),
    .C(_11037_),
    .D(_11043_),
    .X(_11384_));
 sky130_fd_sc_hd__buf_2 _18090_ (.A(_11061_),
    .X(_11385_));
 sky130_fd_sc_hd__buf_2 _18091_ (.A(_11036_),
    .X(_11386_));
 sky130_fd_sc_hd__buf_2 _18092_ (.A(_11057_),
    .X(_11387_));
 sky130_fd_sc_hd__a22oi_1 _18093_ (.A1(_11385_),
    .A2(_11386_),
    .B1(_11157_),
    .B2(_11387_),
    .Y(_11388_));
 sky130_fd_sc_hd__nor2_1 _18094_ (.A(_11384_),
    .B(_11388_),
    .Y(_11389_));
 sky130_fd_sc_hd__xnor2_1 _18095_ (.A(_11383_),
    .B(_11389_),
    .Y(_11390_));
 sky130_fd_sc_hd__o21ba_1 _18096_ (.A1(_11279_),
    .A2(_11283_),
    .B1_N(_11281_),
    .X(_11391_));
 sky130_fd_sc_hd__xnor2_1 _18097_ (.A(_11390_),
    .B(_11391_),
    .Y(_11392_));
 sky130_fd_sc_hd__xnor2_1 _18098_ (.A(_11378_),
    .B(_11392_),
    .Y(_11393_));
 sky130_fd_sc_hd__a21o_1 _18099_ (.A1(_11366_),
    .A2(_11367_),
    .B1(_11393_),
    .X(_11394_));
 sky130_fd_sc_hd__nand3_1 _18100_ (.A(_11366_),
    .B(_11367_),
    .C(_11393_),
    .Y(_11395_));
 sky130_fd_sc_hd__o211ai_2 _18101_ (.A1(_11266_),
    .A2(_11273_),
    .B1(_11394_),
    .C1(_11395_),
    .Y(_11396_));
 sky130_fd_sc_hd__a211o_1 _18102_ (.A1(_11394_),
    .A2(_11395_),
    .B1(_11266_),
    .C1(_11273_),
    .X(_11397_));
 sky130_fd_sc_hd__nand3_1 _18103_ (.A(_11294_),
    .B(_11310_),
    .C(_11311_),
    .Y(_11398_));
 sky130_fd_sc_hd__nand2_1 _18104_ (.A(_11306_),
    .B(_11308_),
    .Y(_11399_));
 sky130_fd_sc_hd__nand2_1 _18105_ (.A(_11300_),
    .B(_11304_),
    .Y(_11400_));
 sky130_fd_sc_hd__a31o_1 _18106_ (.A1(_11245_),
    .A2(_11191_),
    .A3(_11248_),
    .B1(_11247_),
    .X(_11401_));
 sky130_fd_sc_hd__buf_2 _18107_ (.A(_11175_),
    .X(_11402_));
 sky130_fd_sc_hd__nand2_1 _18108_ (.A(_10737_),
    .B(_11402_),
    .Y(_11403_));
 sky130_fd_sc_hd__buf_2 _18109_ (.A(_10912_),
    .X(_11404_));
 sky130_fd_sc_hd__buf_2 _18110_ (.A(_11059_),
    .X(_11405_));
 sky130_fd_sc_hd__nand4_2 _18111_ (.A(_11404_),
    .B(_11299_),
    .C(_11405_),
    .D(_11197_),
    .Y(_11406_));
 sky130_fd_sc_hd__a22o_1 _18112_ (.A1(_11299_),
    .A2(_10973_),
    .B1(_11197_),
    .B2(_11302_),
    .X(_11407_));
 sky130_fd_sc_hd__nand3b_2 _18113_ (.A_N(_11403_),
    .B(_11406_),
    .C(_11407_),
    .Y(_11408_));
 sky130_fd_sc_hd__a21bo_1 _18114_ (.A1(_11406_),
    .A2(_11407_),
    .B1_N(_11403_),
    .X(_11409_));
 sky130_fd_sc_hd__nand3_4 _18115_ (.A(_11401_),
    .B(_11408_),
    .C(_11409_),
    .Y(_11410_));
 sky130_fd_sc_hd__a21o_1 _18116_ (.A1(_11408_),
    .A2(_11409_),
    .B1(_11401_),
    .X(_11411_));
 sky130_fd_sc_hd__nand3_4 _18117_ (.A(_11400_),
    .B(_11410_),
    .C(_11411_),
    .Y(_11412_));
 sky130_fd_sc_hd__a21o_1 _18118_ (.A1(_11410_),
    .A2(_11411_),
    .B1(_11400_),
    .X(_11413_));
 sky130_fd_sc_hd__nand3_4 _18119_ (.A(_11251_),
    .B(_11412_),
    .C(_11413_),
    .Y(_11414_));
 sky130_fd_sc_hd__a21o_1 _18120_ (.A1(_11412_),
    .A2(_11413_),
    .B1(_11251_),
    .X(_11415_));
 sky130_fd_sc_hd__and3_1 _18121_ (.A(_11399_),
    .B(_11414_),
    .C(_11415_),
    .X(_11416_));
 sky130_fd_sc_hd__a21oi_1 _18122_ (.A1(_11414_),
    .A2(_11415_),
    .B1(_11399_),
    .Y(_11417_));
 sky130_fd_sc_hd__a211o_1 _18123_ (.A1(_11310_),
    .A2(_11398_),
    .B1(_11416_),
    .C1(_11417_),
    .X(_11418_));
 sky130_fd_sc_hd__o211ai_2 _18124_ (.A1(_11416_),
    .A2(_11417_),
    .B1(_11310_),
    .C1(_11398_),
    .Y(_11419_));
 sky130_fd_sc_hd__and4_1 _18125_ (.A(_11396_),
    .B(_11397_),
    .C(_11418_),
    .D(_11419_),
    .X(_11420_));
 sky130_fd_sc_hd__a22oi_1 _18126_ (.A1(_11396_),
    .A2(_11397_),
    .B1(_11418_),
    .B2(_11419_),
    .Y(_11421_));
 sky130_fd_sc_hd__a211o_1 _18127_ (.A1(_11364_),
    .A2(_11365_),
    .B1(_11420_),
    .C1(_11421_),
    .X(_11422_));
 sky130_fd_sc_hd__o211ai_1 _18128_ (.A1(_11420_),
    .A2(_11421_),
    .B1(_11364_),
    .C1(_11365_),
    .Y(_11423_));
 sky130_fd_sc_hd__nand3b_1 _18129_ (.A_N(_11363_),
    .B(_11422_),
    .C(_11423_),
    .Y(_11424_));
 sky130_fd_sc_hd__a21bo_1 _18130_ (.A1(_11422_),
    .A2(_11423_),
    .B1_N(_11363_),
    .X(_11425_));
 sky130_fd_sc_hd__nand3b_1 _18131_ (.A_N(_11320_),
    .B(_11424_),
    .C(_11425_),
    .Y(_11426_));
 sky130_fd_sc_hd__a21bo_1 _18132_ (.A1(_11424_),
    .A2(_11425_),
    .B1_N(_11320_),
    .X(_11427_));
 sky130_fd_sc_hd__and3_1 _18133_ (.A(_11342_),
    .B(_11426_),
    .C(_11427_),
    .X(_11428_));
 sky130_fd_sc_hd__a21oi_1 _18134_ (.A1(_11426_),
    .A2(_11427_),
    .B1(_11342_),
    .Y(_11429_));
 sky130_fd_sc_hd__nor2_1 _18135_ (.A(_11428_),
    .B(_11429_),
    .Y(_11430_));
 sky130_fd_sc_hd__nor2_1 _18136_ (.A(_11322_),
    .B(_11328_),
    .Y(_11431_));
 sky130_fd_sc_hd__xnor2_1 _18137_ (.A(_11430_),
    .B(_11431_),
    .Y(_11432_));
 sky130_fd_sc_hd__xor2_1 _18138_ (.A(_11340_),
    .B(_11432_),
    .X(_11433_));
 sky130_fd_sc_hd__or2_1 _18139_ (.A(_11330_),
    .B(_11332_),
    .X(_11434_));
 sky130_fd_sc_hd__xnor2_1 _18140_ (.A(_11433_),
    .B(_11434_),
    .Y(_11435_));
 sky130_fd_sc_hd__o211a_1 _18141_ (.A1(_11332_),
    .A2(_11333_),
    .B1(_11228_),
    .C1(_11229_),
    .X(_11436_));
 sky130_fd_sc_hd__a31oi_1 _18142_ (.A1(_11337_),
    .A2(_11338_),
    .A3(_11334_),
    .B1(_11436_),
    .Y(_11437_));
 sky130_fd_sc_hd__xnor2_1 _18143_ (.A(_11435_),
    .B(_11437_),
    .Y(_00060_));
 sky130_fd_sc_hd__nand2_1 _18144_ (.A(_11433_),
    .B(_11434_),
    .Y(_11438_));
 sky130_fd_sc_hd__a311o_1 _18145_ (.A1(_11337_),
    .A2(_11338_),
    .A3(_11334_),
    .B1(_11436_),
    .C1(_11435_),
    .X(_11439_));
 sky130_fd_sc_hd__and2b_1 _18146_ (.A_N(_11341_),
    .B(_11318_),
    .X(_11440_));
 sky130_fd_sc_hd__nand2_1 _18147_ (.A(_11394_),
    .B(_11396_),
    .Y(_11441_));
 sky130_fd_sc_hd__xnor2_1 _18148_ (.A(_11422_),
    .B(_11441_),
    .Y(_11442_));
 sky130_fd_sc_hd__buf_2 _18149_ (.A(\genblk1.pcpi_mul.rs2[15] ),
    .X(_11443_));
 sky130_fd_sc_hd__clkbuf_4 _18150_ (.A(_11443_),
    .X(_11444_));
 sky130_fd_sc_hd__buf_2 _18151_ (.A(_11444_),
    .X(_11445_));
 sky130_fd_sc_hd__clkbuf_2 _18152_ (.A(_11445_),
    .X(_11446_));
 sky130_fd_sc_hd__buf_4 _18153_ (.A(_11446_),
    .X(_11447_));
 sky130_fd_sc_hd__nand2_1 _18154_ (.A(_10591_),
    .B(_11447_),
    .Y(_11448_));
 sky130_fd_sc_hd__nand2_1 _18155_ (.A(_11404_),
    .B(_10961_),
    .Y(_11449_));
 sky130_fd_sc_hd__and4_1 _18156_ (.A(_10719_),
    .B(_10794_),
    .C(_11141_),
    .D(_11144_),
    .X(_11450_));
 sky130_fd_sc_hd__a22o_1 _18157_ (.A1(_10790_),
    .A2(_10956_),
    .B1(_11107_),
    .B2(_10665_),
    .X(_11451_));
 sky130_fd_sc_hd__and2b_1 _18158_ (.A_N(_11450_),
    .B(_11451_),
    .X(_11452_));
 sky130_fd_sc_hd__xnor2_1 _18159_ (.A(_11449_),
    .B(_11452_),
    .Y(_11453_));
 sky130_fd_sc_hd__nand2_1 _18160_ (.A(_10675_),
    .B(_11350_),
    .Y(_11454_));
 sky130_fd_sc_hd__buf_2 _18161_ (.A(_11352_),
    .X(_11455_));
 sky130_fd_sc_hd__and4_1 _18162_ (.A(_10634_),
    .B(_10628_),
    .C(_11235_),
    .D(_11455_),
    .X(_11456_));
 sky130_fd_sc_hd__clkbuf_2 _18163_ (.A(\genblk1.pcpi_mul.rs2[14] ),
    .X(_11457_));
 sky130_fd_sc_hd__clkbuf_4 _18164_ (.A(_11457_),
    .X(_11458_));
 sky130_fd_sc_hd__a22oi_2 _18165_ (.A1(_10607_),
    .A2(_11356_),
    .B1(_11458_),
    .B2(_10786_),
    .Y(_11459_));
 sky130_fd_sc_hd__or3_1 _18166_ (.A(_11454_),
    .B(_11456_),
    .C(_11459_),
    .X(_11460_));
 sky130_fd_sc_hd__o21ai_1 _18167_ (.A1(_11456_),
    .A2(_11459_),
    .B1(_11454_),
    .Y(_11461_));
 sky130_fd_sc_hd__a21bo_1 _18168_ (.A1(_11351_),
    .A2(_11357_),
    .B1_N(_11355_),
    .X(_11462_));
 sky130_fd_sc_hd__and3_1 _18169_ (.A(_11460_),
    .B(_11461_),
    .C(_11462_),
    .X(_11463_));
 sky130_fd_sc_hd__a21o_1 _18170_ (.A1(_11460_),
    .A2(_11461_),
    .B1(_11462_),
    .X(_11464_));
 sky130_fd_sc_hd__and2b_1 _18171_ (.A_N(_11463_),
    .B(_11464_),
    .X(_11465_));
 sky130_fd_sc_hd__xnor2_1 _18172_ (.A(_11453_),
    .B(_11465_),
    .Y(_11466_));
 sky130_fd_sc_hd__or2_1 _18173_ (.A(_11448_),
    .B(_11466_),
    .X(_11467_));
 sky130_fd_sc_hd__nand2_1 _18174_ (.A(_11448_),
    .B(_11466_),
    .Y(_11468_));
 sky130_fd_sc_hd__and2_1 _18175_ (.A(_11467_),
    .B(_11468_),
    .X(_11469_));
 sky130_fd_sc_hd__nand4_1 _18176_ (.A(_11396_),
    .B(_11397_),
    .C(_11418_),
    .D(_11419_),
    .Y(_11470_));
 sky130_fd_sc_hd__or2b_1 _18177_ (.A(_11391_),
    .B_N(_11390_),
    .X(_11471_));
 sky130_fd_sc_hd__nand2_1 _18178_ (.A(_11378_),
    .B(_11392_),
    .Y(_11472_));
 sky130_fd_sc_hd__clkbuf_2 _18179_ (.A(_11171_),
    .X(_11473_));
 sky130_fd_sc_hd__clkbuf_4 _18180_ (.A(_11473_),
    .X(_11474_));
 sky130_fd_sc_hd__nand2_1 _18181_ (.A(_10633_),
    .B(_11369_),
    .Y(_11475_));
 sky130_fd_sc_hd__buf_2 _18182_ (.A(_11379_),
    .X(_11476_));
 sky130_fd_sc_hd__buf_2 _18183_ (.A(_11476_),
    .X(_11477_));
 sky130_fd_sc_hd__nand2_1 _18184_ (.A(_10641_),
    .B(_11477_),
    .Y(_11478_));
 sky130_fd_sc_hd__buf_2 _18185_ (.A(_11372_),
    .X(_11479_));
 sky130_fd_sc_hd__clkbuf_2 _18186_ (.A(\genblk1.pcpi_mul.rs1[14] ),
    .X(_11480_));
 sky130_fd_sc_hd__buf_2 _18187_ (.A(_11480_),
    .X(_11481_));
 sky130_fd_sc_hd__clkbuf_4 _18188_ (.A(_11481_),
    .X(_11482_));
 sky130_fd_sc_hd__and4_2 _18189_ (.A(_11044_),
    .B(_10632_),
    .C(_11479_),
    .D(_11482_),
    .X(_11483_));
 sky130_fd_sc_hd__a21oi_1 _18190_ (.A1(_11475_),
    .A2(_11478_),
    .B1(_11483_),
    .Y(_11484_));
 sky130_fd_sc_hd__a21oi_1 _18191_ (.A1(_10680_),
    .A2(_11474_),
    .B1(_11484_),
    .Y(_11485_));
 sky130_fd_sc_hd__and3_1 _18192_ (.A(_10626_),
    .B(_11474_),
    .C(_11484_),
    .X(_11486_));
 sky130_fd_sc_hd__nor2_1 _18193_ (.A(_11485_),
    .B(_11486_),
    .Y(_11487_));
 sky130_fd_sc_hd__clkbuf_2 _18194_ (.A(\genblk1.pcpi_mul.rs1[15] ),
    .X(_11488_));
 sky130_fd_sc_hd__clkbuf_4 _18195_ (.A(_11488_),
    .X(_11489_));
 sky130_fd_sc_hd__clkbuf_2 _18196_ (.A(_11489_),
    .X(_11490_));
 sky130_fd_sc_hd__buf_2 _18197_ (.A(_11490_),
    .X(_11491_));
 sky130_fd_sc_hd__nand2_1 _18198_ (.A(_11053_),
    .B(_11491_),
    .Y(_11492_));
 sky130_fd_sc_hd__and4_1 _18199_ (.A(_10662_),
    .B(_11058_),
    .C(_11156_),
    .D(_11160_),
    .X(_11493_));
 sky130_fd_sc_hd__a22oi_1 _18200_ (.A1(_11282_),
    .A2(_11039_),
    .B1(_11056_),
    .B2(_10672_),
    .Y(_11494_));
 sky130_fd_sc_hd__nor2_1 _18201_ (.A(_11493_),
    .B(_11494_),
    .Y(_11495_));
 sky130_fd_sc_hd__xnor2_1 _18202_ (.A(_11492_),
    .B(_11495_),
    .Y(_11496_));
 sky130_fd_sc_hd__o21ba_1 _18203_ (.A1(_11383_),
    .A2(_11388_),
    .B1_N(_11384_),
    .X(_11497_));
 sky130_fd_sc_hd__xnor2_1 _18204_ (.A(_11496_),
    .B(_11497_),
    .Y(_11498_));
 sky130_fd_sc_hd__xnor2_1 _18205_ (.A(_11487_),
    .B(_11498_),
    .Y(_11499_));
 sky130_fd_sc_hd__a21o_1 _18206_ (.A1(_11471_),
    .A2(_11472_),
    .B1(_11499_),
    .X(_11500_));
 sky130_fd_sc_hd__nand3_1 _18207_ (.A(_11471_),
    .B(_11472_),
    .C(_11499_),
    .Y(_11501_));
 sky130_fd_sc_hd__o211a_1 _18208_ (.A1(_11374_),
    .A2(_11377_),
    .B1(_11500_),
    .C1(_11501_),
    .X(_11502_));
 sky130_fd_sc_hd__a211oi_1 _18209_ (.A1(_11500_),
    .A2(_11501_),
    .B1(_11374_),
    .C1(_11377_),
    .Y(_11503_));
 sky130_fd_sc_hd__nand3_2 _18210_ (.A(_11399_),
    .B(_11414_),
    .C(_11415_),
    .Y(_11504_));
 sky130_fd_sc_hd__a21o_1 _18211_ (.A1(_11348_),
    .A2(_11361_),
    .B1(_11360_),
    .X(_11505_));
 sky130_fd_sc_hd__nand2_1 _18212_ (.A(_11406_),
    .B(_11408_),
    .Y(_11506_));
 sky130_fd_sc_hd__a31o_1 _18213_ (.A1(_11343_),
    .A2(_11191_),
    .A3(_11346_),
    .B1(_11345_),
    .X(_11507_));
 sky130_fd_sc_hd__clkbuf_4 _18214_ (.A(_10787_),
    .X(_11508_));
 sky130_fd_sc_hd__nand2_1 _18215_ (.A(_11508_),
    .B(_11042_),
    .Y(_11509_));
 sky130_fd_sc_hd__nand4_2 _18216_ (.A(_10783_),
    .B(_10973_),
    .C(_11201_),
    .D(_11177_),
    .Y(_11510_));
 sky130_fd_sc_hd__a22o_1 _18217_ (.A1(_11059_),
    .A2(_11201_),
    .B1(_11177_),
    .B2(_11084_),
    .X(_11511_));
 sky130_fd_sc_hd__nand3b_1 _18218_ (.A_N(_11509_),
    .B(_11510_),
    .C(_11511_),
    .Y(_11512_));
 sky130_fd_sc_hd__a21bo_1 _18219_ (.A1(_11510_),
    .A2(_11511_),
    .B1_N(_11509_),
    .X(_11513_));
 sky130_fd_sc_hd__nand3_2 _18220_ (.A(_11507_),
    .B(_11512_),
    .C(_11513_),
    .Y(_11514_));
 sky130_fd_sc_hd__a21o_1 _18221_ (.A1(_11512_),
    .A2(_11513_),
    .B1(_11507_),
    .X(_11515_));
 sky130_fd_sc_hd__nand3_2 _18222_ (.A(_11506_),
    .B(_11514_),
    .C(_11515_),
    .Y(_11516_));
 sky130_fd_sc_hd__a21o_1 _18223_ (.A1(_11514_),
    .A2(_11515_),
    .B1(_11506_),
    .X(_11517_));
 sky130_fd_sc_hd__and3_2 _18224_ (.A(_11505_),
    .B(_11516_),
    .C(_11517_),
    .X(_11518_));
 sky130_fd_sc_hd__a21oi_2 _18225_ (.A1(_11516_),
    .A2(_11517_),
    .B1(_11505_),
    .Y(_11519_));
 sky130_fd_sc_hd__a211oi_4 _18226_ (.A1(_11410_),
    .A2(_11412_),
    .B1(_11518_),
    .C1(_11519_),
    .Y(_11520_));
 sky130_fd_sc_hd__o211a_1 _18227_ (.A1(_11518_),
    .A2(_11519_),
    .B1(_11410_),
    .C1(_11412_),
    .X(_11521_));
 sky130_fd_sc_hd__a211oi_4 _18228_ (.A1(_11414_),
    .A2(_11504_),
    .B1(_11520_),
    .C1(_11521_),
    .Y(_11522_));
 sky130_fd_sc_hd__o211a_1 _18229_ (.A1(_11520_),
    .A2(_11521_),
    .B1(_11414_),
    .C1(_11504_),
    .X(_11523_));
 sky130_fd_sc_hd__nor4_1 _18230_ (.A(_11502_),
    .B(_11503_),
    .C(_11522_),
    .D(_11523_),
    .Y(_11524_));
 sky130_fd_sc_hd__o22a_1 _18231_ (.A1(_11502_),
    .A2(_11503_),
    .B1(_11522_),
    .B2(_11523_),
    .X(_11525_));
 sky130_fd_sc_hd__a211o_1 _18232_ (.A1(_11418_),
    .A2(_11470_),
    .B1(net352),
    .C1(_11525_),
    .X(_11526_));
 sky130_fd_sc_hd__o211ai_1 _18233_ (.A1(net352),
    .A2(_11525_),
    .B1(_11418_),
    .C1(_11470_),
    .Y(_11527_));
 sky130_fd_sc_hd__and3_1 _18234_ (.A(_11469_),
    .B(_11526_),
    .C(_11527_),
    .X(_11528_));
 sky130_fd_sc_hd__a21oi_1 _18235_ (.A1(_11526_),
    .A2(_11527_),
    .B1(_11469_),
    .Y(_11529_));
 sky130_fd_sc_hd__or3_1 _18236_ (.A(_11424_),
    .B(_11528_),
    .C(_11529_),
    .X(_11530_));
 sky130_fd_sc_hd__o21ai_1 _18237_ (.A1(_11528_),
    .A2(_11529_),
    .B1(_11424_),
    .Y(_11531_));
 sky130_fd_sc_hd__nand3_1 _18238_ (.A(_11442_),
    .B(_11530_),
    .C(_11531_),
    .Y(_11532_));
 sky130_fd_sc_hd__a21o_1 _18239_ (.A1(_11530_),
    .A2(_11531_),
    .B1(_11442_),
    .X(_11533_));
 sky130_fd_sc_hd__a21bo_1 _18240_ (.A1(_11342_),
    .A2(_11427_),
    .B1_N(_11426_),
    .X(_11534_));
 sky130_fd_sc_hd__nand3_1 _18241_ (.A(_11532_),
    .B(_11533_),
    .C(_11534_),
    .Y(_11535_));
 sky130_fd_sc_hd__a21o_1 _18242_ (.A1(_11532_),
    .A2(_11533_),
    .B1(_11534_),
    .X(_11536_));
 sky130_fd_sc_hd__and3_1 _18243_ (.A(_11440_),
    .B(_11535_),
    .C(_11536_),
    .X(_11537_));
 sky130_fd_sc_hd__a21oi_1 _18244_ (.A1(_11535_),
    .A2(_11536_),
    .B1(_11440_),
    .Y(_11538_));
 sky130_fd_sc_hd__or2_1 _18245_ (.A(_11537_),
    .B(_11538_),
    .X(_11539_));
 sky130_fd_sc_hd__or3_1 _18246_ (.A(_11428_),
    .B(_11429_),
    .C(_11431_),
    .X(_11540_));
 sky130_fd_sc_hd__a21boi_1 _18247_ (.A1(_11340_),
    .A2(_11432_),
    .B1_N(_11540_),
    .Y(_11541_));
 sky130_fd_sc_hd__or2_1 _18248_ (.A(_11539_),
    .B(_11541_),
    .X(_11542_));
 sky130_fd_sc_hd__nand2_1 _18249_ (.A(_11539_),
    .B(_11541_),
    .Y(_11543_));
 sky130_fd_sc_hd__nand2_1 _18250_ (.A(_11542_),
    .B(_11543_),
    .Y(_11544_));
 sky130_fd_sc_hd__a21oi_1 _18251_ (.A1(_11438_),
    .A2(_11439_),
    .B1(_11544_),
    .Y(_11545_));
 sky130_fd_sc_hd__and3_1 _18252_ (.A(_11438_),
    .B(_11439_),
    .C(_11544_),
    .X(_11546_));
 sky130_fd_sc_hd__nor2_1 _18253_ (.A(_11545_),
    .B(_11546_),
    .Y(_00061_));
 sky130_fd_sc_hd__a21o_1 _18254_ (.A1(_11438_),
    .A2(_11439_),
    .B1(_11544_),
    .X(_11547_));
 sky130_fd_sc_hd__and2_1 _18255_ (.A(_11542_),
    .B(_11547_),
    .X(_11548_));
 sky130_vsdinv _18256_ (.A(_11537_),
    .Y(_11549_));
 sky130_fd_sc_hd__or2b_1 _18257_ (.A(_11422_),
    .B_N(_11441_),
    .X(_11550_));
 sky130_fd_sc_hd__a21oi_1 _18258_ (.A1(_11471_),
    .A2(_11472_),
    .B1(_11499_),
    .Y(_11551_));
 sky130_fd_sc_hd__or2_1 _18259_ (.A(_11551_),
    .B(_11502_),
    .X(_11552_));
 sky130_fd_sc_hd__xor2_1 _18260_ (.A(_11526_),
    .B(_11552_),
    .X(_11553_));
 sky130_fd_sc_hd__buf_2 _18261_ (.A(\genblk1.pcpi_mul.rs2[16] ),
    .X(_11554_));
 sky130_fd_sc_hd__buf_2 _18262_ (.A(_11554_),
    .X(_11555_));
 sky130_fd_sc_hd__clkbuf_2 _18263_ (.A(_11555_),
    .X(_11556_));
 sky130_fd_sc_hd__clkbuf_4 _18264_ (.A(_11556_),
    .X(_11557_));
 sky130_fd_sc_hd__a22oi_1 _18265_ (.A1(_10597_),
    .A2(_11447_),
    .B1(_11557_),
    .B2(_10591_),
    .Y(_11558_));
 sky130_fd_sc_hd__buf_2 _18266_ (.A(_11443_),
    .X(_11559_));
 sky130_fd_sc_hd__clkbuf_4 _18267_ (.A(_11559_),
    .X(_11560_));
 sky130_fd_sc_hd__clkbuf_2 _18268_ (.A(_11560_),
    .X(_11561_));
 sky130_fd_sc_hd__and4_2 _18269_ (.A(_10623_),
    .B(_10596_),
    .C(_11561_),
    .D(_11557_),
    .X(_11562_));
 sky130_fd_sc_hd__nand2_1 _18270_ (.A(_11405_),
    .B(_10961_),
    .Y(_11563_));
 sky130_fd_sc_hd__and4_1 _18271_ (.A(_11301_),
    .B(_10794_),
    .C(_11141_),
    .D(_11144_),
    .X(_11564_));
 sky130_fd_sc_hd__a22o_1 _18272_ (.A1(_11301_),
    .A2(_10956_),
    .B1(_11107_),
    .B2(_10790_),
    .X(_11565_));
 sky130_fd_sc_hd__and2b_1 _18273_ (.A_N(_11564_),
    .B(_11565_),
    .X(_11566_));
 sky130_fd_sc_hd__xnor2_1 _18274_ (.A(_11563_),
    .B(_11566_),
    .Y(_11567_));
 sky130_fd_sc_hd__nand2_1 _18275_ (.A(_10744_),
    .B(_11350_),
    .Y(_11568_));
 sky130_fd_sc_hd__and4_1 _18276_ (.A(_10628_),
    .B(_10861_),
    .C(_11235_),
    .D(_11455_),
    .X(_11569_));
 sky130_fd_sc_hd__a22oi_2 _18277_ (.A1(_10717_),
    .A2(_11356_),
    .B1(_11458_),
    .B2(_10607_),
    .Y(_11570_));
 sky130_fd_sc_hd__or3_1 _18278_ (.A(_11568_),
    .B(_11569_),
    .C(_11570_),
    .X(_11571_));
 sky130_fd_sc_hd__o21ai_1 _18279_ (.A1(_11569_),
    .A2(_11570_),
    .B1(_11568_),
    .Y(_11572_));
 sky130_fd_sc_hd__o21bai_1 _18280_ (.A1(_11454_),
    .A2(_11459_),
    .B1_N(_11456_),
    .Y(_11573_));
 sky130_fd_sc_hd__and3_1 _18281_ (.A(_11571_),
    .B(_11572_),
    .C(_11573_),
    .X(_11574_));
 sky130_fd_sc_hd__a21o_1 _18282_ (.A1(_11571_),
    .A2(_11572_),
    .B1(_11573_),
    .X(_11575_));
 sky130_fd_sc_hd__and2b_1 _18283_ (.A_N(_11574_),
    .B(_11575_),
    .X(_11576_));
 sky130_fd_sc_hd__xnor2_1 _18284_ (.A(_11567_),
    .B(_11576_),
    .Y(_11577_));
 sky130_fd_sc_hd__nor3_1 _18285_ (.A(_11558_),
    .B(_11562_),
    .C(_11577_),
    .Y(_11578_));
 sky130_fd_sc_hd__o21a_1 _18286_ (.A1(_11558_),
    .A2(_11562_),
    .B1(_11577_),
    .X(_11579_));
 sky130_fd_sc_hd__or2_1 _18287_ (.A(_11578_),
    .B(_11579_),
    .X(_11580_));
 sky130_fd_sc_hd__or2_1 _18288_ (.A(_11467_),
    .B(_11580_),
    .X(_11581_));
 sky130_fd_sc_hd__nand2_1 _18289_ (.A(_11467_),
    .B(_11580_),
    .Y(_11582_));
 sky130_fd_sc_hd__and2_1 _18290_ (.A(_11581_),
    .B(_11582_),
    .X(_11583_));
 sky130_fd_sc_hd__or2b_1 _18291_ (.A(_11497_),
    .B_N(_11496_),
    .X(_11584_));
 sky130_fd_sc_hd__nand2_1 _18292_ (.A(_11487_),
    .B(_11498_),
    .Y(_11585_));
 sky130_fd_sc_hd__nand2_1 _18293_ (.A(_10633_),
    .B(_11382_),
    .Y(_11586_));
 sky130_fd_sc_hd__nand2_2 _18294_ (.A(_10600_),
    .B(_11490_),
    .Y(_11587_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18295_ (.A(\genblk1.pcpi_mul.rs1[15] ),
    .X(_11588_));
 sky130_fd_sc_hd__clkbuf_2 _18296_ (.A(_11588_),
    .X(_11589_));
 sky130_fd_sc_hd__buf_4 _18297_ (.A(_11589_),
    .X(_11590_));
 sky130_fd_sc_hd__buf_2 _18298_ (.A(_11590_),
    .X(_11591_));
 sky130_fd_sc_hd__nand2_2 _18299_ (.A(_10632_),
    .B(_11591_),
    .Y(_11592_));
 sky130_fd_sc_hd__nor2_1 _18300_ (.A(_11478_),
    .B(_11592_),
    .Y(_11593_));
 sky130_fd_sc_hd__a21oi_1 _18301_ (.A1(_11586_),
    .A2(_11587_),
    .B1(_11593_),
    .Y(_11594_));
 sky130_fd_sc_hd__nand2_1 _18302_ (.A(_10626_),
    .B(_11369_),
    .Y(_11595_));
 sky130_fd_sc_hd__xnor2_1 _18303_ (.A(_11594_),
    .B(_11595_),
    .Y(_11596_));
 sky130_fd_sc_hd__clkbuf_2 _18304_ (.A(\genblk1.pcpi_mul.rs1[16] ),
    .X(_11597_));
 sky130_fd_sc_hd__clkbuf_4 _18305_ (.A(_11597_),
    .X(_11598_));
 sky130_fd_sc_hd__clkbuf_4 _18306_ (.A(_11598_),
    .X(_11599_));
 sky130_fd_sc_hd__nand2_1 _18307_ (.A(_11053_),
    .B(_11599_),
    .Y(_11600_));
 sky130_fd_sc_hd__clkbuf_2 _18308_ (.A(_11170_),
    .X(_11601_));
 sky130_fd_sc_hd__and4_1 _18309_ (.A(_11063_),
    .B(_11061_),
    .C(_11055_),
    .D(_11601_),
    .X(_11602_));
 sky130_fd_sc_hd__a22oi_1 _18310_ (.A1(_11058_),
    .A2(_11160_),
    .B1(_11265_),
    .B2(_10662_),
    .Y(_11603_));
 sky130_fd_sc_hd__nor2_1 _18311_ (.A(_11602_),
    .B(_11603_),
    .Y(_11604_));
 sky130_fd_sc_hd__xnor2_2 _18312_ (.A(_11600_),
    .B(_11604_),
    .Y(_11605_));
 sky130_fd_sc_hd__o21ba_1 _18313_ (.A1(_11492_),
    .A2(_11494_),
    .B1_N(_11493_),
    .X(_11606_));
 sky130_fd_sc_hd__xnor2_1 _18314_ (.A(_11605_),
    .B(_11606_),
    .Y(_11607_));
 sky130_fd_sc_hd__xnor2_1 _18315_ (.A(_11596_),
    .B(_11607_),
    .Y(_11608_));
 sky130_fd_sc_hd__a21o_1 _18316_ (.A1(_11584_),
    .A2(_11585_),
    .B1(_11608_),
    .X(_11609_));
 sky130_fd_sc_hd__nand3_2 _18317_ (.A(_11584_),
    .B(_11585_),
    .C(_11608_),
    .Y(_11610_));
 sky130_fd_sc_hd__o211ai_4 _18318_ (.A1(_11483_),
    .A2(_11486_),
    .B1(_11609_),
    .C1(_11610_),
    .Y(_11611_));
 sky130_fd_sc_hd__a211o_1 _18319_ (.A1(_11609_),
    .A2(_11610_),
    .B1(_11483_),
    .C1(_11486_),
    .X(_11612_));
 sky130_fd_sc_hd__a21o_1 _18320_ (.A1(_11453_),
    .A2(_11464_),
    .B1(_11463_),
    .X(_11613_));
 sky130_fd_sc_hd__nand2_1 _18321_ (.A(_11510_),
    .B(_11512_),
    .Y(_11614_));
 sky130_fd_sc_hd__a31o_1 _18322_ (.A1(_11193_),
    .A2(_11190_),
    .A3(_11451_),
    .B1(_11450_),
    .X(_11615_));
 sky130_fd_sc_hd__nand2_1 _18323_ (.A(_10736_),
    .B(_11269_),
    .Y(_11616_));
 sky130_fd_sc_hd__nand4_2 _18324_ (.A(_11298_),
    .B(_11196_),
    .C(_11048_),
    .D(_11036_),
    .Y(_11617_));
 sky130_fd_sc_hd__a22o_1 _18325_ (.A1(_10998_),
    .A2(_10967_),
    .B1(_10969_),
    .B2(_11082_),
    .X(_11618_));
 sky130_fd_sc_hd__nand3b_1 _18326_ (.A_N(_11616_),
    .B(_11617_),
    .C(_11618_),
    .Y(_11619_));
 sky130_fd_sc_hd__a21bo_1 _18327_ (.A1(_11617_),
    .A2(_11618_),
    .B1_N(_11616_),
    .X(_11620_));
 sky130_fd_sc_hd__nand3_2 _18328_ (.A(_11615_),
    .B(_11619_),
    .C(_11620_),
    .Y(_11621_));
 sky130_fd_sc_hd__a21o_1 _18329_ (.A1(_11619_),
    .A2(_11620_),
    .B1(_11615_),
    .X(_11622_));
 sky130_fd_sc_hd__nand3_2 _18330_ (.A(_11614_),
    .B(_11621_),
    .C(_11622_),
    .Y(_11623_));
 sky130_fd_sc_hd__a21o_1 _18331_ (.A1(_11621_),
    .A2(_11622_),
    .B1(_11614_),
    .X(_11624_));
 sky130_fd_sc_hd__and3_1 _18332_ (.A(_11613_),
    .B(_11623_),
    .C(_11624_),
    .X(_11625_));
 sky130_fd_sc_hd__a21oi_1 _18333_ (.A1(_11623_),
    .A2(_11624_),
    .B1(_11613_),
    .Y(_11626_));
 sky130_fd_sc_hd__a211o_2 _18334_ (.A1(_11514_),
    .A2(_11516_),
    .B1(_11625_),
    .C1(_11626_),
    .X(_11627_));
 sky130_fd_sc_hd__o211ai_2 _18335_ (.A1(_11625_),
    .A2(_11626_),
    .B1(_11514_),
    .C1(_11516_),
    .Y(_11628_));
 sky130_fd_sc_hd__o211ai_4 _18336_ (.A1(_11518_),
    .A2(_11520_),
    .B1(_11627_),
    .C1(_11628_),
    .Y(_11629_));
 sky130_fd_sc_hd__a211o_1 _18337_ (.A1(_11627_),
    .A2(_11628_),
    .B1(_11518_),
    .C1(_11520_),
    .X(_11630_));
 sky130_fd_sc_hd__nand4_4 _18338_ (.A(_11611_),
    .B(_11612_),
    .C(_11629_),
    .D(_11630_),
    .Y(_11631_));
 sky130_fd_sc_hd__a22o_1 _18339_ (.A1(_11611_),
    .A2(_11612_),
    .B1(_11629_),
    .B2(_11630_),
    .X(_11632_));
 sky130_fd_sc_hd__o211ai_4 _18340_ (.A1(_11522_),
    .A2(net351),
    .B1(_11631_),
    .C1(_11632_),
    .Y(_11633_));
 sky130_fd_sc_hd__a211o_1 _18341_ (.A1(_11631_),
    .A2(_11632_),
    .B1(_11522_),
    .C1(net352),
    .X(_11634_));
 sky130_fd_sc_hd__and3_1 _18342_ (.A(_11583_),
    .B(_11633_),
    .C(_11634_),
    .X(_11635_));
 sky130_fd_sc_hd__a21o_1 _18343_ (.A1(_11633_),
    .A2(_11634_),
    .B1(_11583_),
    .X(_11636_));
 sky130_fd_sc_hd__or2b_1 _18344_ (.A(_11635_),
    .B_N(_11636_),
    .X(_11637_));
 sky130_fd_sc_hd__xnor2_1 _18345_ (.A(_11528_),
    .B(_11637_),
    .Y(_11638_));
 sky130_fd_sc_hd__xnor2_1 _18346_ (.A(_11553_),
    .B(_11638_),
    .Y(_11639_));
 sky130_fd_sc_hd__nand2_1 _18347_ (.A(_11530_),
    .B(_11532_),
    .Y(_11640_));
 sky130_fd_sc_hd__xnor2_1 _18348_ (.A(_11639_),
    .B(_11640_),
    .Y(_11641_));
 sky130_fd_sc_hd__xnor2_1 _18349_ (.A(_11550_),
    .B(_11641_),
    .Y(_11642_));
 sky130_fd_sc_hd__a21oi_1 _18350_ (.A1(_11535_),
    .A2(_11549_),
    .B1(_11642_),
    .Y(_11643_));
 sky130_fd_sc_hd__and3_1 _18351_ (.A(_11535_),
    .B(_11549_),
    .C(_11642_),
    .X(_11644_));
 sky130_fd_sc_hd__or2_1 _18352_ (.A(_11643_),
    .B(_11644_),
    .X(_11645_));
 sky130_fd_sc_hd__nor2_1 _18353_ (.A(_11548_),
    .B(_11645_),
    .Y(_11646_));
 sky130_fd_sc_hd__and3_1 _18354_ (.A(_11542_),
    .B(_11547_),
    .C(_11645_),
    .X(_11647_));
 sky130_fd_sc_hd__nor2_1 _18355_ (.A(_11646_),
    .B(_11647_),
    .Y(_00062_));
 sky130_fd_sc_hd__and2_1 _18356_ (.A(_11639_),
    .B(_11640_),
    .X(_11648_));
 sky130_fd_sc_hd__nor2_1 _18357_ (.A(_11550_),
    .B(_11641_),
    .Y(_11649_));
 sky130_fd_sc_hd__or2b_1 _18358_ (.A(_11526_),
    .B_N(_11552_),
    .X(_11650_));
 sky130_fd_sc_hd__and3b_1 _18359_ (.A_N(_11635_),
    .B(_11636_),
    .C(_11528_),
    .X(_11651_));
 sky130_fd_sc_hd__and2b_1 _18360_ (.A_N(_11553_),
    .B(_11638_),
    .X(_11652_));
 sky130_fd_sc_hd__nand2_1 _18361_ (.A(_11609_),
    .B(_11611_),
    .Y(_11653_));
 sky130_fd_sc_hd__xor2_1 _18362_ (.A(_11633_),
    .B(_11653_),
    .X(_11654_));
 sky130_fd_sc_hd__nand2_1 _18363_ (.A(_10609_),
    .B(_11445_),
    .Y(_11655_));
 sky130_fd_sc_hd__clkbuf_2 _18364_ (.A(_11555_),
    .X(_11656_));
 sky130_fd_sc_hd__clkbuf_2 _18365_ (.A(\genblk1.pcpi_mul.rs2[17] ),
    .X(_11657_));
 sky130_fd_sc_hd__buf_2 _18366_ (.A(_11657_),
    .X(_11658_));
 sky130_fd_sc_hd__clkbuf_2 _18367_ (.A(_11658_),
    .X(_11659_));
 sky130_fd_sc_hd__and4_1 _18368_ (.A(_11113_),
    .B(_10638_),
    .C(_11656_),
    .D(_11659_),
    .X(_11660_));
 sky130_fd_sc_hd__clkbuf_2 _18369_ (.A(\genblk1.pcpi_mul.rs2[16] ),
    .X(_11661_));
 sky130_fd_sc_hd__buf_2 _18370_ (.A(_11661_),
    .X(_11662_));
 sky130_fd_sc_hd__buf_2 _18371_ (.A(_11662_),
    .X(_11663_));
 sky130_fd_sc_hd__clkbuf_4 _18372_ (.A(_11663_),
    .X(_11664_));
 sky130_fd_sc_hd__clkbuf_2 _18373_ (.A(_11658_),
    .X(_11665_));
 sky130_fd_sc_hd__buf_4 _18374_ (.A(_11665_),
    .X(_11666_));
 sky130_fd_sc_hd__a22oi_4 _18375_ (.A1(_10636_),
    .A2(_11664_),
    .B1(_11666_),
    .B2(_11113_),
    .Y(_11667_));
 sky130_fd_sc_hd__nor2_1 _18376_ (.A(_11660_),
    .B(_11667_),
    .Y(_11668_));
 sky130_fd_sc_hd__xnor2_1 _18377_ (.A(_11655_),
    .B(_11668_),
    .Y(_11669_));
 sky130_fd_sc_hd__and2_1 _18378_ (.A(_11562_),
    .B(_11669_),
    .X(_11670_));
 sky130_fd_sc_hd__nor2_1 _18379_ (.A(_11562_),
    .B(_11669_),
    .Y(_11671_));
 sky130_fd_sc_hd__or2_1 _18380_ (.A(_11670_),
    .B(_11671_),
    .X(_11672_));
 sky130_fd_sc_hd__nand2_1 _18381_ (.A(_11402_),
    .B(_10893_),
    .Y(_11673_));
 sky130_fd_sc_hd__and4_1 _18382_ (.A(_11301_),
    .B(_10852_),
    .C(_10956_),
    .D(_11107_),
    .X(_11674_));
 sky130_fd_sc_hd__a22o_1 _18383_ (.A1(_10852_),
    .A2(_10956_),
    .B1(_11107_),
    .B2(_11301_),
    .X(_11675_));
 sky130_fd_sc_hd__and2b_1 _18384_ (.A_N(_11674_),
    .B(_11675_),
    .X(_11676_));
 sky130_fd_sc_hd__xnor2_2 _18385_ (.A(_11673_),
    .B(_11676_),
    .Y(_11677_));
 sky130_fd_sc_hd__nand2_1 _18386_ (.A(_10746_),
    .B(_11350_),
    .Y(_11678_));
 sky130_fd_sc_hd__and4_1 _18387_ (.A(_10861_),
    .B(_10719_),
    .C(_11356_),
    .D(_11458_),
    .X(_11679_));
 sky130_fd_sc_hd__a22oi_2 _18388_ (.A1(_10665_),
    .A2(_11356_),
    .B1(_11354_),
    .B2(_10675_),
    .Y(_11680_));
 sky130_fd_sc_hd__or3_1 _18389_ (.A(_11678_),
    .B(_11679_),
    .C(_11680_),
    .X(_11681_));
 sky130_fd_sc_hd__o21ai_1 _18390_ (.A1(_11679_),
    .A2(_11680_),
    .B1(_11678_),
    .Y(_11682_));
 sky130_fd_sc_hd__o21bai_1 _18391_ (.A1(_11568_),
    .A2(_11570_),
    .B1_N(_11569_),
    .Y(_11683_));
 sky130_fd_sc_hd__and3_1 _18392_ (.A(_11681_),
    .B(_11682_),
    .C(_11683_),
    .X(_11684_));
 sky130_fd_sc_hd__a21o_1 _18393_ (.A1(_11681_),
    .A2(_11682_),
    .B1(_11683_),
    .X(_11685_));
 sky130_fd_sc_hd__and2b_1 _18394_ (.A_N(_11684_),
    .B(_11685_),
    .X(_11686_));
 sky130_fd_sc_hd__xnor2_1 _18395_ (.A(_11677_),
    .B(_11686_),
    .Y(_11687_));
 sky130_fd_sc_hd__or2_1 _18396_ (.A(_11672_),
    .B(_11687_),
    .X(_11688_));
 sky130_fd_sc_hd__nand2_1 _18397_ (.A(_11672_),
    .B(_11687_),
    .Y(_11689_));
 sky130_fd_sc_hd__and3_1 _18398_ (.A(_11578_),
    .B(_11688_),
    .C(_11689_),
    .X(_11690_));
 sky130_fd_sc_hd__a21oi_1 _18399_ (.A1(_11688_),
    .A2(_11689_),
    .B1(_11578_),
    .Y(_11691_));
 sky130_fd_sc_hd__nand2_1 _18400_ (.A(_11629_),
    .B(_11631_),
    .Y(_11692_));
 sky130_fd_sc_hd__or2_1 _18401_ (.A(_11478_),
    .B(_11592_),
    .X(_11693_));
 sky130_fd_sc_hd__a211o_1 _18402_ (.A1(_11586_),
    .A2(_11587_),
    .B1(_11593_),
    .C1(_11595_),
    .X(_11694_));
 sky130_fd_sc_hd__or2b_1 _18403_ (.A(_11606_),
    .B_N(_11605_),
    .X(_11695_));
 sky130_fd_sc_hd__nand2_1 _18404_ (.A(_11596_),
    .B(_11607_),
    .Y(_11696_));
 sky130_fd_sc_hd__buf_1 _18405_ (.A(\genblk1.pcpi_mul.rs1[16] ),
    .X(_11697_));
 sky130_fd_sc_hd__buf_2 _18406_ (.A(_11697_),
    .X(_11698_));
 sky130_fd_sc_hd__clkbuf_4 _18407_ (.A(_11698_),
    .X(_11699_));
 sky130_fd_sc_hd__nand2_2 _18408_ (.A(_11044_),
    .B(_11699_),
    .Y(_11700_));
 sky130_fd_sc_hd__nand2_1 _18409_ (.A(_11041_),
    .B(_11699_),
    .Y(_11701_));
 sky130_fd_sc_hd__nor2_1 _18410_ (.A(_11587_),
    .B(_11701_),
    .Y(_11702_));
 sky130_fd_sc_hd__a21oi_1 _18411_ (.A1(_11592_),
    .A2(_11700_),
    .B1(_11702_),
    .Y(_11703_));
 sky130_fd_sc_hd__buf_2 _18412_ (.A(_10644_),
    .X(_11704_));
 sky130_fd_sc_hd__nand2_1 _18413_ (.A(_11704_),
    .B(_11382_),
    .Y(_11705_));
 sky130_fd_sc_hd__xnor2_1 _18414_ (.A(_11703_),
    .B(_11705_),
    .Y(_11706_));
 sky130_fd_sc_hd__buf_2 _18415_ (.A(\genblk1.pcpi_mul.rs1[17] ),
    .X(_11707_));
 sky130_fd_sc_hd__buf_4 _18416_ (.A(_11707_),
    .X(_11708_));
 sky130_fd_sc_hd__nand2_1 _18417_ (.A(_10669_),
    .B(_11708_),
    .Y(_11709_));
 sky130_fd_sc_hd__buf_2 _18418_ (.A(_10699_),
    .X(_11710_));
 sky130_fd_sc_hd__buf_2 _18419_ (.A(_10701_),
    .X(_11711_));
 sky130_fd_sc_hd__buf_2 _18420_ (.A(_11371_),
    .X(_11712_));
 sky130_fd_sc_hd__and4_1 _18421_ (.A(_11710_),
    .B(_11711_),
    .C(_11171_),
    .D(_11712_),
    .X(_11713_));
 sky130_fd_sc_hd__a22oi_1 _18422_ (.A1(_11061_),
    .A2(_11601_),
    .B1(_11277_),
    .B2(_11057_),
    .Y(_11714_));
 sky130_fd_sc_hd__nor2_1 _18423_ (.A(_11713_),
    .B(_11714_),
    .Y(_11715_));
 sky130_fd_sc_hd__xnor2_2 _18424_ (.A(_11709_),
    .B(_11715_),
    .Y(_11716_));
 sky130_fd_sc_hd__o21ba_1 _18425_ (.A1(_11600_),
    .A2(_11603_),
    .B1_N(_11602_),
    .X(_11717_));
 sky130_fd_sc_hd__xnor2_1 _18426_ (.A(_11716_),
    .B(_11717_),
    .Y(_11718_));
 sky130_fd_sc_hd__xnor2_1 _18427_ (.A(_11706_),
    .B(_11718_),
    .Y(_11719_));
 sky130_fd_sc_hd__a21oi_1 _18428_ (.A1(_11695_),
    .A2(_11696_),
    .B1(_11719_),
    .Y(_11720_));
 sky130_fd_sc_hd__and3_1 _18429_ (.A(_11695_),
    .B(_11696_),
    .C(_11719_),
    .X(_11721_));
 sky130_fd_sc_hd__a211oi_2 _18430_ (.A1(_11693_),
    .A2(_11694_),
    .B1(_11720_),
    .C1(_11721_),
    .Y(_11722_));
 sky130_fd_sc_hd__o211a_1 _18431_ (.A1(_11720_),
    .A2(_11721_),
    .B1(_11693_),
    .C1(_11694_),
    .X(_11723_));
 sky130_fd_sc_hd__nand3_1 _18432_ (.A(_11613_),
    .B(_11623_),
    .C(_11624_),
    .Y(_11724_));
 sky130_fd_sc_hd__a21o_1 _18433_ (.A1(_11567_),
    .A2(_11575_),
    .B1(_11574_),
    .X(_11725_));
 sky130_fd_sc_hd__nand2_1 _18434_ (.A(_11617_),
    .B(_11619_),
    .Y(_11726_));
 sky130_fd_sc_hd__a31o_1 _18435_ (.A1(_10973_),
    .A2(_11190_),
    .A3(_11565_),
    .B1(_11564_),
    .X(_11727_));
 sky130_fd_sc_hd__buf_2 _18436_ (.A(_11159_),
    .X(_11728_));
 sky130_fd_sc_hd__nand4_2 _18437_ (.A(_11298_),
    .B(_11196_),
    .C(_11036_),
    .D(_11038_),
    .Y(_11729_));
 sky130_fd_sc_hd__a22o_1 _18438_ (.A1(_10998_),
    .A2(_10969_),
    .B1(_11155_),
    .B2(_11082_),
    .X(_11730_));
 sky130_fd_sc_hd__nand4_2 _18439_ (.A(_11089_),
    .B(_11728_),
    .C(_11729_),
    .D(_11730_),
    .Y(_11731_));
 sky130_fd_sc_hd__a22o_1 _18440_ (.A1(_11508_),
    .A2(_11264_),
    .B1(_11729_),
    .B2(_11730_),
    .X(_11732_));
 sky130_fd_sc_hd__nand3_2 _18441_ (.A(_11727_),
    .B(_11731_),
    .C(_11732_),
    .Y(_11733_));
 sky130_fd_sc_hd__a21o_1 _18442_ (.A1(_11731_),
    .A2(_11732_),
    .B1(_11727_),
    .X(_11734_));
 sky130_fd_sc_hd__nand3_2 _18443_ (.A(_11726_),
    .B(_11733_),
    .C(_11734_),
    .Y(_11735_));
 sky130_fd_sc_hd__a21o_1 _18444_ (.A1(_11733_),
    .A2(_11734_),
    .B1(_11726_),
    .X(_11736_));
 sky130_fd_sc_hd__and3_2 _18445_ (.A(_11725_),
    .B(_11735_),
    .C(_11736_),
    .X(_11737_));
 sky130_fd_sc_hd__a21oi_2 _18446_ (.A1(_11735_),
    .A2(_11736_),
    .B1(_11725_),
    .Y(_11738_));
 sky130_fd_sc_hd__a211oi_4 _18447_ (.A1(_11621_),
    .A2(_11623_),
    .B1(_11737_),
    .C1(_11738_),
    .Y(_11739_));
 sky130_fd_sc_hd__o211a_1 _18448_ (.A1(_11737_),
    .A2(_11738_),
    .B1(_11621_),
    .C1(_11623_),
    .X(_11740_));
 sky130_fd_sc_hd__a211oi_2 _18449_ (.A1(_11724_),
    .A2(_11627_),
    .B1(_11739_),
    .C1(_11740_),
    .Y(_11741_));
 sky130_fd_sc_hd__o211a_1 _18450_ (.A1(_11739_),
    .A2(_11740_),
    .B1(_11724_),
    .C1(_11627_),
    .X(_11742_));
 sky130_fd_sc_hd__nor4_1 _18451_ (.A(_11722_),
    .B(_11723_),
    .C(_11741_),
    .D(_11742_),
    .Y(_11743_));
 sky130_fd_sc_hd__o22a_1 _18452_ (.A1(_11722_),
    .A2(_11723_),
    .B1(_11741_),
    .B2(_11742_),
    .X(_11744_));
 sky130_fd_sc_hd__or3_1 _18453_ (.A(_11581_),
    .B(net350),
    .C(_11744_),
    .X(_11745_));
 sky130_fd_sc_hd__o21ai_1 _18454_ (.A1(net350),
    .A2(_11744_),
    .B1(_11581_),
    .Y(_11746_));
 sky130_fd_sc_hd__nand3_1 _18455_ (.A(_11692_),
    .B(_11745_),
    .C(_11746_),
    .Y(_11747_));
 sky130_fd_sc_hd__a21o_1 _18456_ (.A1(_11745_),
    .A2(_11746_),
    .B1(_11692_),
    .X(_11748_));
 sky130_fd_sc_hd__or4bb_1 _18457_ (.A(_11690_),
    .B(_11691_),
    .C_N(_11747_),
    .D_N(_11748_),
    .X(_11749_));
 sky130_fd_sc_hd__a2bb2o_1 _18458_ (.A1_N(_11690_),
    .A2_N(_11691_),
    .B1(_11747_),
    .B2(_11748_),
    .X(_11750_));
 sky130_fd_sc_hd__and3_1 _18459_ (.A(_11635_),
    .B(_11749_),
    .C(_11750_),
    .X(_11751_));
 sky130_fd_sc_hd__a21oi_1 _18460_ (.A1(_11749_),
    .A2(_11750_),
    .B1(_11635_),
    .Y(_11752_));
 sky130_fd_sc_hd__or3_2 _18461_ (.A(_11654_),
    .B(_11751_),
    .C(_11752_),
    .X(_11753_));
 sky130_fd_sc_hd__o21ai_1 _18462_ (.A1(_11751_),
    .A2(_11752_),
    .B1(_11654_),
    .Y(_11754_));
 sky130_fd_sc_hd__o211a_1 _18463_ (.A1(_11651_),
    .A2(_11652_),
    .B1(_11753_),
    .C1(_11754_),
    .X(_11755_));
 sky130_fd_sc_hd__a211oi_1 _18464_ (.A1(_11753_),
    .A2(_11754_),
    .B1(_11651_),
    .C1(_11652_),
    .Y(_11756_));
 sky130_fd_sc_hd__or3_1 _18465_ (.A(_11650_),
    .B(_11755_),
    .C(_11756_),
    .X(_11757_));
 sky130_fd_sc_hd__o21ai_1 _18466_ (.A1(_11755_),
    .A2(_11756_),
    .B1(_11650_),
    .Y(_11758_));
 sky130_fd_sc_hd__o211a_1 _18467_ (.A1(_11648_),
    .A2(_11649_),
    .B1(_11757_),
    .C1(_11758_),
    .X(_11759_));
 sky130_fd_sc_hd__a211oi_1 _18468_ (.A1(_11757_),
    .A2(_11758_),
    .B1(_11648_),
    .C1(_11649_),
    .Y(_11760_));
 sky130_fd_sc_hd__nor2_1 _18469_ (.A(_11759_),
    .B(_11760_),
    .Y(_11761_));
 sky130_fd_sc_hd__nor2_1 _18470_ (.A(_11643_),
    .B(_11646_),
    .Y(_11762_));
 sky130_fd_sc_hd__xnor2_1 _18471_ (.A(_11761_),
    .B(_11762_),
    .Y(_00063_));
 sky130_vsdinv _18472_ (.A(_11755_),
    .Y(_11763_));
 sky130_fd_sc_hd__or2b_1 _18473_ (.A(_11633_),
    .B_N(_11653_),
    .X(_11764_));
 sky130_vsdinv _18474_ (.A(_11751_),
    .Y(_11765_));
 sky130_fd_sc_hd__nand2_1 _18475_ (.A(_11745_),
    .B(_11747_),
    .Y(_11766_));
 sky130_fd_sc_hd__nor2_1 _18476_ (.A(_11720_),
    .B(_11722_),
    .Y(_11767_));
 sky130_fd_sc_hd__xnor2_1 _18477_ (.A(_11766_),
    .B(_11767_),
    .Y(_11768_));
 sky130_fd_sc_hd__clkbuf_2 _18478_ (.A(\genblk1.pcpi_mul.rs2[18] ),
    .X(_11769_));
 sky130_fd_sc_hd__buf_2 _18479_ (.A(_11769_),
    .X(_11770_));
 sky130_fd_sc_hd__buf_2 _18480_ (.A(_11770_),
    .X(_11771_));
 sky130_fd_sc_hd__clkbuf_4 _18481_ (.A(_11771_),
    .X(_11772_));
 sky130_fd_sc_hd__buf_4 _18482_ (.A(_11772_),
    .X(_11773_));
 sky130_fd_sc_hd__nand2_1 _18483_ (.A(_10603_),
    .B(_11773_),
    .Y(_11774_));
 sky130_fd_sc_hd__buf_2 _18484_ (.A(_11559_),
    .X(_11775_));
 sky130_fd_sc_hd__nand2_2 _18485_ (.A(_10651_),
    .B(_11775_),
    .Y(_11776_));
 sky130_fd_sc_hd__buf_2 _18486_ (.A(_10752_),
    .X(_11777_));
 sky130_fd_sc_hd__buf_2 _18487_ (.A(_11777_),
    .X(_11778_));
 sky130_fd_sc_hd__and4_1 _18488_ (.A(_10595_),
    .B(_11778_),
    .C(_11556_),
    .D(_11659_),
    .X(_11779_));
 sky130_fd_sc_hd__clkbuf_2 _18489_ (.A(\genblk1.pcpi_mul.rs2[17] ),
    .X(_11780_));
 sky130_fd_sc_hd__buf_2 _18490_ (.A(_11780_),
    .X(_11781_));
 sky130_fd_sc_hd__clkbuf_4 _18491_ (.A(_11781_),
    .X(_11782_));
 sky130_fd_sc_hd__a22oi_2 _18492_ (.A1(_10608_),
    .A2(_11664_),
    .B1(_11782_),
    .B2(_10636_),
    .Y(_11783_));
 sky130_fd_sc_hd__nor2_2 _18493_ (.A(_11779_),
    .B(_11783_),
    .Y(_11784_));
 sky130_fd_sc_hd__xnor2_4 _18494_ (.A(_11776_),
    .B(_11784_),
    .Y(_11785_));
 sky130_fd_sc_hd__o21ba_1 _18495_ (.A1(_11655_),
    .A2(_11667_),
    .B1_N(_11660_),
    .X(_11786_));
 sky130_fd_sc_hd__xnor2_1 _18496_ (.A(_11785_),
    .B(_11786_),
    .Y(_11787_));
 sky130_fd_sc_hd__xnor2_1 _18497_ (.A(_11670_),
    .B(_11787_),
    .Y(_11788_));
 sky130_fd_sc_hd__nand2_1 _18498_ (.A(_10893_),
    .B(_11386_),
    .Y(_11789_));
 sky130_fd_sc_hd__and4_1 _18499_ (.A(_11062_),
    .B(_11048_),
    .C(_10963_),
    .D(_11111_),
    .X(_11790_));
 sky130_fd_sc_hd__a22o_1 _18500_ (.A1(_11048_),
    .A2(_10963_),
    .B1(_11111_),
    .B2(_11062_),
    .X(_11791_));
 sky130_fd_sc_hd__and2b_1 _18501_ (.A_N(_11790_),
    .B(_11791_),
    .X(_11792_));
 sky130_fd_sc_hd__xnor2_2 _18502_ (.A(_11789_),
    .B(_11792_),
    .Y(_11793_));
 sky130_fd_sc_hd__nand2_1 _18503_ (.A(_10912_),
    .B(_11350_),
    .Y(_11794_));
 sky130_fd_sc_hd__clkbuf_4 _18504_ (.A(\genblk1.pcpi_mul.rs2[13] ),
    .X(_11795_));
 sky130_fd_sc_hd__and4_1 _18505_ (.A(_10741_),
    .B(_10745_),
    .C(_11795_),
    .D(_11353_),
    .X(_11796_));
 sky130_fd_sc_hd__a22oi_2 _18506_ (.A1(_10746_),
    .A2(_11241_),
    .B1(_11354_),
    .B2(_10744_),
    .Y(_11797_));
 sky130_fd_sc_hd__or3_1 _18507_ (.A(_11794_),
    .B(_11796_),
    .C(_11797_),
    .X(_11798_));
 sky130_fd_sc_hd__o21ai_1 _18508_ (.A1(_11796_),
    .A2(_11797_),
    .B1(_11794_),
    .Y(_11799_));
 sky130_fd_sc_hd__o21bai_1 _18509_ (.A1(_11678_),
    .A2(_11680_),
    .B1_N(_11679_),
    .Y(_11800_));
 sky130_fd_sc_hd__and3_1 _18510_ (.A(_11798_),
    .B(_11799_),
    .C(_11800_),
    .X(_11801_));
 sky130_fd_sc_hd__a21o_1 _18511_ (.A1(_11798_),
    .A2(_11799_),
    .B1(_11800_),
    .X(_11802_));
 sky130_fd_sc_hd__and2b_1 _18512_ (.A_N(_11801_),
    .B(_11802_),
    .X(_11803_));
 sky130_fd_sc_hd__xnor2_1 _18513_ (.A(_11793_),
    .B(_11803_),
    .Y(_11804_));
 sky130_fd_sc_hd__nor2_1 _18514_ (.A(_11788_),
    .B(_11804_),
    .Y(_11805_));
 sky130_fd_sc_hd__and2_1 _18515_ (.A(_11788_),
    .B(_11804_),
    .X(_11806_));
 sky130_fd_sc_hd__or3_1 _18516_ (.A(_11688_),
    .B(_11805_),
    .C(_11806_),
    .X(_11807_));
 sky130_fd_sc_hd__o21ai_1 _18517_ (.A1(_11805_),
    .A2(_11806_),
    .B1(_11688_),
    .Y(_11808_));
 sky130_fd_sc_hd__nand2_1 _18518_ (.A(_11807_),
    .B(_11808_),
    .Y(_11809_));
 sky130_fd_sc_hd__or2_1 _18519_ (.A(_11774_),
    .B(_11809_),
    .X(_11810_));
 sky130_fd_sc_hd__nand2_1 _18520_ (.A(_11774_),
    .B(_11809_),
    .Y(_11811_));
 sky130_fd_sc_hd__and2_1 _18521_ (.A(_11810_),
    .B(_11811_),
    .X(_11812_));
 sky130_fd_sc_hd__nor2_1 _18522_ (.A(_11741_),
    .B(_11743_),
    .Y(_11813_));
 sky130_fd_sc_hd__or2_1 _18523_ (.A(_11587_),
    .B(_11701_),
    .X(_11814_));
 sky130_fd_sc_hd__a211o_1 _18524_ (.A1(_11592_),
    .A2(_11700_),
    .B1(_11702_),
    .C1(_11705_),
    .X(_11815_));
 sky130_fd_sc_hd__or2b_1 _18525_ (.A(_11717_),
    .B_N(_11716_),
    .X(_11816_));
 sky130_fd_sc_hd__nand2_1 _18526_ (.A(_11706_),
    .B(_11718_),
    .Y(_11817_));
 sky130_fd_sc_hd__clkbuf_2 _18527_ (.A(\genblk1.pcpi_mul.rs1[17] ),
    .X(_11818_));
 sky130_fd_sc_hd__clkbuf_4 _18528_ (.A(_11818_),
    .X(_11819_));
 sky130_fd_sc_hd__buf_2 _18529_ (.A(_11819_),
    .X(_11820_));
 sky130_fd_sc_hd__nand2_2 _18530_ (.A(_10641_),
    .B(_11820_),
    .Y(_11821_));
 sky130_fd_sc_hd__nand2_2 _18531_ (.A(_11041_),
    .B(_11708_),
    .Y(_11822_));
 sky130_fd_sc_hd__nor2_1 _18532_ (.A(_11700_),
    .B(_11822_),
    .Y(_11823_));
 sky130_fd_sc_hd__a21oi_1 _18533_ (.A1(_11701_),
    .A2(_11821_),
    .B1(_11823_),
    .Y(_11824_));
 sky130_fd_sc_hd__clkbuf_4 _18534_ (.A(_11589_),
    .X(_11825_));
 sky130_fd_sc_hd__buf_4 _18535_ (.A(_11825_),
    .X(_11826_));
 sky130_fd_sc_hd__nand2_1 _18536_ (.A(_11704_),
    .B(_11826_),
    .Y(_11827_));
 sky130_fd_sc_hd__xnor2_1 _18537_ (.A(_11824_),
    .B(_11827_),
    .Y(_11828_));
 sky130_fd_sc_hd__clkbuf_2 _18538_ (.A(\genblk1.pcpi_mul.rs1[18] ),
    .X(_11829_));
 sky130_fd_sc_hd__clkbuf_4 _18539_ (.A(_11829_),
    .X(_11830_));
 sky130_fd_sc_hd__clkbuf_4 _18540_ (.A(_11830_),
    .X(_11831_));
 sky130_fd_sc_hd__nand2_1 _18541_ (.A(_10669_),
    .B(_11831_),
    .Y(_11832_));
 sky130_fd_sc_hd__and4_1 _18542_ (.A(_10671_),
    .B(_11711_),
    .C(_11712_),
    .D(_11476_),
    .X(_11833_));
 sky130_fd_sc_hd__clkbuf_4 _18543_ (.A(_11481_),
    .X(_11834_));
 sky130_fd_sc_hd__a22oi_1 _18544_ (.A1(_11061_),
    .A2(_11372_),
    .B1(_11834_),
    .B2(_11057_),
    .Y(_11835_));
 sky130_fd_sc_hd__nor2_1 _18545_ (.A(_11833_),
    .B(_11835_),
    .Y(_11836_));
 sky130_fd_sc_hd__xnor2_2 _18546_ (.A(_11832_),
    .B(_11836_),
    .Y(_11837_));
 sky130_fd_sc_hd__o21ba_1 _18547_ (.A1(_11709_),
    .A2(_11714_),
    .B1_N(_11713_),
    .X(_11838_));
 sky130_fd_sc_hd__xnor2_1 _18548_ (.A(_11837_),
    .B(_11838_),
    .Y(_11839_));
 sky130_fd_sc_hd__xnor2_1 _18549_ (.A(_11828_),
    .B(_11839_),
    .Y(_11840_));
 sky130_fd_sc_hd__a21oi_1 _18550_ (.A1(_11816_),
    .A2(_11817_),
    .B1(_11840_),
    .Y(_11841_));
 sky130_fd_sc_hd__and3_1 _18551_ (.A(_11816_),
    .B(_11817_),
    .C(_11840_),
    .X(_11842_));
 sky130_fd_sc_hd__a211oi_1 _18552_ (.A1(_11814_),
    .A2(_11815_),
    .B1(_11841_),
    .C1(_11842_),
    .Y(_11843_));
 sky130_fd_sc_hd__o211a_1 _18553_ (.A1(_11841_),
    .A2(_11842_),
    .B1(_11814_),
    .C1(_11815_),
    .X(_11844_));
 sky130_fd_sc_hd__a21o_1 _18554_ (.A1(_11677_),
    .A2(_11685_),
    .B1(_11684_),
    .X(_11845_));
 sky130_fd_sc_hd__nand2_1 _18555_ (.A(_11729_),
    .B(_11731_),
    .Y(_11846_));
 sky130_fd_sc_hd__a31o_1 _18556_ (.A1(_11049_),
    .A2(_11190_),
    .A3(_11675_),
    .B1(_11674_),
    .X(_11847_));
 sky130_fd_sc_hd__nand2_1 _18557_ (.A(_11508_),
    .B(_11261_),
    .Y(_11848_));
 sky130_fd_sc_hd__nand4_2 _18558_ (.A(_11084_),
    .B(_11086_),
    .C(_11038_),
    .D(_11055_),
    .Y(_11849_));
 sky130_fd_sc_hd__a22o_1 _18559_ (.A1(_11196_),
    .A2(_11155_),
    .B1(_11067_),
    .B2(_11298_),
    .X(_11850_));
 sky130_fd_sc_hd__nand3b_1 _18560_ (.A_N(_11848_),
    .B(_11849_),
    .C(_11850_),
    .Y(_11851_));
 sky130_fd_sc_hd__a21bo_1 _18561_ (.A1(_11849_),
    .A2(_11850_),
    .B1_N(_11848_),
    .X(_11852_));
 sky130_fd_sc_hd__nand3_2 _18562_ (.A(_11847_),
    .B(_11851_),
    .C(_11852_),
    .Y(_11853_));
 sky130_fd_sc_hd__a21o_1 _18563_ (.A1(_11851_),
    .A2(_11852_),
    .B1(_11847_),
    .X(_11854_));
 sky130_fd_sc_hd__nand3_2 _18564_ (.A(_11846_),
    .B(_11853_),
    .C(_11854_),
    .Y(_11855_));
 sky130_fd_sc_hd__a21o_1 _18565_ (.A1(_11853_),
    .A2(_11854_),
    .B1(_11846_),
    .X(_11856_));
 sky130_fd_sc_hd__and3_1 _18566_ (.A(_11845_),
    .B(_11855_),
    .C(_11856_),
    .X(_11857_));
 sky130_fd_sc_hd__a21oi_1 _18567_ (.A1(_11855_),
    .A2(_11856_),
    .B1(_11845_),
    .Y(_11858_));
 sky130_fd_sc_hd__a211o_2 _18568_ (.A1(_11733_),
    .A2(_11735_),
    .B1(_11857_),
    .C1(_11858_),
    .X(_11859_));
 sky130_fd_sc_hd__o211ai_2 _18569_ (.A1(_11857_),
    .A2(_11858_),
    .B1(_11733_),
    .C1(_11735_),
    .Y(_11860_));
 sky130_fd_sc_hd__o211ai_4 _18570_ (.A1(_11737_),
    .A2(_11739_),
    .B1(_11859_),
    .C1(_11860_),
    .Y(_11861_));
 sky130_fd_sc_hd__a211o_1 _18571_ (.A1(_11859_),
    .A2(_11860_),
    .B1(_11737_),
    .C1(_11739_),
    .X(_11862_));
 sky130_fd_sc_hd__or4bb_2 _18572_ (.A(_11843_),
    .B(_11844_),
    .C_N(_11861_),
    .D_N(_11862_),
    .X(_11863_));
 sky130_fd_sc_hd__a2bb2o_1 _18573_ (.A1_N(_11843_),
    .A2_N(_11844_),
    .B1(_11861_),
    .B2(_11862_),
    .X(_11864_));
 sky130_fd_sc_hd__and3_1 _18574_ (.A(_11690_),
    .B(_11863_),
    .C(_11864_),
    .X(_11865_));
 sky130_fd_sc_hd__a21oi_1 _18575_ (.A1(_11863_),
    .A2(_11864_),
    .B1(_11690_),
    .Y(_11866_));
 sky130_fd_sc_hd__or3_1 _18576_ (.A(_11813_),
    .B(_11865_),
    .C(_11866_),
    .X(_11867_));
 sky130_fd_sc_hd__o21ai_1 _18577_ (.A1(_11865_),
    .A2(_11866_),
    .B1(_11813_),
    .Y(_11868_));
 sky130_fd_sc_hd__and3_1 _18578_ (.A(_11812_),
    .B(_11867_),
    .C(_11868_),
    .X(_11869_));
 sky130_fd_sc_hd__a21oi_1 _18579_ (.A1(_11867_),
    .A2(_11868_),
    .B1(_11812_),
    .Y(_11870_));
 sky130_fd_sc_hd__or3_2 _18580_ (.A(_11749_),
    .B(_11869_),
    .C(_11870_),
    .X(_11871_));
 sky130_fd_sc_hd__o21ai_1 _18581_ (.A1(_11869_),
    .A2(_11870_),
    .B1(_11749_),
    .Y(_11872_));
 sky130_fd_sc_hd__and3_1 _18582_ (.A(_11768_),
    .B(_11871_),
    .C(_11872_),
    .X(_11873_));
 sky130_fd_sc_hd__a21oi_1 _18583_ (.A1(_11871_),
    .A2(_11872_),
    .B1(_11768_),
    .Y(_11874_));
 sky130_fd_sc_hd__a211oi_2 _18584_ (.A1(_11765_),
    .A2(_11753_),
    .B1(_11873_),
    .C1(_11874_),
    .Y(_11875_));
 sky130_fd_sc_hd__o211a_1 _18585_ (.A1(_11873_),
    .A2(_11874_),
    .B1(_11765_),
    .C1(_11753_),
    .X(_11876_));
 sky130_fd_sc_hd__nor3_1 _18586_ (.A(_11764_),
    .B(_11875_),
    .C(_11876_),
    .Y(_11877_));
 sky130_fd_sc_hd__o21a_1 _18587_ (.A1(_11875_),
    .A2(_11876_),
    .B1(_11764_),
    .X(_11878_));
 sky130_fd_sc_hd__a211oi_1 _18588_ (.A1(_11763_),
    .A2(_11757_),
    .B1(_11877_),
    .C1(_11878_),
    .Y(_11879_));
 sky130_fd_sc_hd__o211a_1 _18589_ (.A1(_11877_),
    .A2(_11878_),
    .B1(_11763_),
    .C1(_11757_),
    .X(_11880_));
 sky130_fd_sc_hd__nor2_1 _18590_ (.A(_11879_),
    .B(_11880_),
    .Y(_11881_));
 sky130_fd_sc_hd__o21ba_1 _18591_ (.A1(_11643_),
    .A2(_11759_),
    .B1_N(_11760_),
    .X(_11882_));
 sky130_fd_sc_hd__a21o_1 _18592_ (.A1(_11646_),
    .A2(_11761_),
    .B1(_11882_),
    .X(_11883_));
 sky130_fd_sc_hd__xor2_1 _18593_ (.A(_11881_),
    .B(_11883_),
    .X(_00064_));
 sky130_fd_sc_hd__a21o_1 _18594_ (.A1(_11745_),
    .A2(_11747_),
    .B1(_11767_),
    .X(_11884_));
 sky130_fd_sc_hd__nand3_1 _18595_ (.A(_11768_),
    .B(_11871_),
    .C(_11872_),
    .Y(_11885_));
 sky130_fd_sc_hd__and2b_1 _18596_ (.A_N(_11865_),
    .B(_11867_),
    .X(_11886_));
 sky130_fd_sc_hd__nor2_1 _18597_ (.A(_11841_),
    .B(_11843_),
    .Y(_11887_));
 sky130_fd_sc_hd__xnor2_1 _18598_ (.A(_11886_),
    .B(_11887_),
    .Y(_11888_));
 sky130_fd_sc_hd__clkbuf_2 _18599_ (.A(\genblk1.pcpi_mul.rs2[19] ),
    .X(_11889_));
 sky130_fd_sc_hd__buf_2 _18600_ (.A(_11889_),
    .X(_11890_));
 sky130_fd_sc_hd__clkbuf_4 _18601_ (.A(_11890_),
    .X(_11891_));
 sky130_fd_sc_hd__buf_4 _18602_ (.A(_11891_),
    .X(_11892_));
 sky130_fd_sc_hd__a22oi_4 _18603_ (.A1(_10598_),
    .A2(_11773_),
    .B1(_11892_),
    .B2(_10592_),
    .Y(_11893_));
 sky130_fd_sc_hd__clkbuf_2 _18604_ (.A(\genblk1.pcpi_mul.rs2[18] ),
    .X(_11894_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18605_ (.A(_11894_),
    .X(_11895_));
 sky130_fd_sc_hd__buf_2 _18606_ (.A(_11890_),
    .X(_11896_));
 sky130_fd_sc_hd__and4_2 _18607_ (.A(_11113_),
    .B(_10638_),
    .C(_11895_),
    .D(_11896_),
    .X(_11897_));
 sky130_fd_sc_hd__nor2_1 _18608_ (.A(_11893_),
    .B(_11897_),
    .Y(_11898_));
 sky130_fd_sc_hd__and2_1 _18609_ (.A(_11670_),
    .B(_11787_),
    .X(_11899_));
 sky130_fd_sc_hd__clkbuf_4 _18610_ (.A(\genblk1.pcpi_mul.rs2[9] ),
    .X(_11900_));
 sky130_fd_sc_hd__nand2_1 _18611_ (.A(_11900_),
    .B(_11156_),
    .Y(_11901_));
 sky130_fd_sc_hd__and4_1 _18612_ (.A(_11047_),
    .B(_10968_),
    .C(_10962_),
    .D(_11110_),
    .X(_11902_));
 sky130_fd_sc_hd__buf_2 _18613_ (.A(\genblk1.pcpi_mul.rs1[9] ),
    .X(_11903_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18614_ (.A(_11140_),
    .X(_11904_));
 sky130_fd_sc_hd__clkbuf_2 _18615_ (.A(_11143_),
    .X(_11905_));
 sky130_fd_sc_hd__a22o_1 _18616_ (.A1(_11903_),
    .A2(_11904_),
    .B1(_11905_),
    .B2(_11047_),
    .X(_11906_));
 sky130_fd_sc_hd__and2b_1 _18617_ (.A_N(_11902_),
    .B(_11906_),
    .X(_11907_));
 sky130_fd_sc_hd__xnor2_1 _18618_ (.A(_11901_),
    .B(_11907_),
    .Y(_11908_));
 sky130_fd_sc_hd__nand2_1 _18619_ (.A(_10805_),
    .B(_11134_),
    .Y(_11909_));
 sky130_fd_sc_hd__clkbuf_2 _18620_ (.A(_11352_),
    .X(_11910_));
 sky130_fd_sc_hd__and4_1 _18621_ (.A(_10978_),
    .B(_10793_),
    .C(_11240_),
    .D(_11910_),
    .X(_11911_));
 sky130_fd_sc_hd__a22oi_2 _18622_ (.A1(_10848_),
    .A2(_11235_),
    .B1(_11455_),
    .B2(_10696_),
    .Y(_11912_));
 sky130_fd_sc_hd__or3_1 _18623_ (.A(_11909_),
    .B(_11911_),
    .C(_11912_),
    .X(_11913_));
 sky130_fd_sc_hd__o21ai_1 _18624_ (.A1(_11911_),
    .A2(_11912_),
    .B1(_11909_),
    .Y(_11914_));
 sky130_fd_sc_hd__o21bai_1 _18625_ (.A1(_11794_),
    .A2(_11797_),
    .B1_N(_11796_),
    .Y(_11915_));
 sky130_fd_sc_hd__and3_1 _18626_ (.A(_11913_),
    .B(_11914_),
    .C(_11915_),
    .X(_11916_));
 sky130_fd_sc_hd__a21o_1 _18627_ (.A1(_11913_),
    .A2(_11914_),
    .B1(_11915_),
    .X(_11917_));
 sky130_fd_sc_hd__and2b_1 _18628_ (.A_N(_11916_),
    .B(_11917_),
    .X(_11918_));
 sky130_fd_sc_hd__xnor2_1 _18629_ (.A(_11908_),
    .B(_11918_),
    .Y(_11919_));
 sky130_fd_sc_hd__and2b_1 _18630_ (.A_N(_11786_),
    .B(_11785_),
    .X(_11920_));
 sky130_fd_sc_hd__nand2_2 _18631_ (.A(_11245_),
    .B(_11445_),
    .Y(_11921_));
 sky130_fd_sc_hd__clkbuf_2 _18632_ (.A(\genblk1.pcpi_mul.rs2[16] ),
    .X(_11922_));
 sky130_fd_sc_hd__buf_2 _18633_ (.A(_11922_),
    .X(_11923_));
 sky130_fd_sc_hd__buf_2 _18634_ (.A(\genblk1.pcpi_mul.rs2[17] ),
    .X(_11924_));
 sky130_fd_sc_hd__buf_2 _18635_ (.A(_11924_),
    .X(_11925_));
 sky130_fd_sc_hd__and4_1 _18636_ (.A(_10629_),
    .B(_11087_),
    .C(_11923_),
    .D(_11925_),
    .X(_11926_));
 sky130_fd_sc_hd__clkbuf_2 _18637_ (.A(_11781_),
    .X(_11927_));
 sky130_fd_sc_hd__a22oi_1 _18638_ (.A1(_10650_),
    .A2(_11656_),
    .B1(_11927_),
    .B2(_11778_),
    .Y(_11928_));
 sky130_fd_sc_hd__nor2_2 _18639_ (.A(_11926_),
    .B(_11928_),
    .Y(_11929_));
 sky130_fd_sc_hd__xnor2_4 _18640_ (.A(_11921_),
    .B(_11929_),
    .Y(_11930_));
 sky130_fd_sc_hd__o21ba_2 _18641_ (.A1(_11776_),
    .A2(_11783_),
    .B1_N(_11779_),
    .X(_11931_));
 sky130_fd_sc_hd__xnor2_1 _18642_ (.A(_11930_),
    .B(_11931_),
    .Y(_11932_));
 sky130_fd_sc_hd__xnor2_1 _18643_ (.A(_11920_),
    .B(_11932_),
    .Y(_11933_));
 sky130_fd_sc_hd__or2_2 _18644_ (.A(_11919_),
    .B(_11933_),
    .X(_11934_));
 sky130_fd_sc_hd__nand2_1 _18645_ (.A(_11919_),
    .B(_11933_),
    .Y(_11935_));
 sky130_fd_sc_hd__o211a_1 _18646_ (.A1(_11899_),
    .A2(_11805_),
    .B1(_11934_),
    .C1(_11935_),
    .X(_11936_));
 sky130_fd_sc_hd__a211oi_1 _18647_ (.A1(_11934_),
    .A2(_11935_),
    .B1(_11899_),
    .C1(_11805_),
    .Y(_11937_));
 sky130_fd_sc_hd__nor2_1 _18648_ (.A(_11936_),
    .B(_11937_),
    .Y(_11938_));
 sky130_fd_sc_hd__xnor2_1 _18649_ (.A(_11898_),
    .B(_11938_),
    .Y(_11939_));
 sky130_fd_sc_hd__xor2_1 _18650_ (.A(_11810_),
    .B(_11939_),
    .X(_11940_));
 sky130_fd_sc_hd__or2_1 _18651_ (.A(_11700_),
    .B(_11822_),
    .X(_11941_));
 sky130_fd_sc_hd__a211o_1 _18652_ (.A1(_11701_),
    .A2(_11821_),
    .B1(_11823_),
    .C1(_11827_),
    .X(_11942_));
 sky130_fd_sc_hd__or2b_1 _18653_ (.A(_11838_),
    .B_N(_11837_),
    .X(_11943_));
 sky130_fd_sc_hd__nand2_1 _18654_ (.A(_11828_),
    .B(_11839_),
    .Y(_11944_));
 sky130_fd_sc_hd__clkbuf_2 _18655_ (.A(\genblk1.pcpi_mul.rs1[18] ),
    .X(_11945_));
 sky130_fd_sc_hd__clkbuf_4 _18656_ (.A(_11945_),
    .X(_11946_));
 sky130_fd_sc_hd__clkbuf_4 _18657_ (.A(_11946_),
    .X(_11947_));
 sky130_fd_sc_hd__nand2_4 _18658_ (.A(_10600_),
    .B(_11947_),
    .Y(_11948_));
 sky130_fd_sc_hd__clkbuf_4 _18659_ (.A(_11829_),
    .X(_11949_));
 sky130_fd_sc_hd__clkbuf_4 _18660_ (.A(_11949_),
    .X(_11950_));
 sky130_fd_sc_hd__nand2_2 _18661_ (.A(_10632_),
    .B(_11950_),
    .Y(_11951_));
 sky130_fd_sc_hd__nor2_1 _18662_ (.A(_11821_),
    .B(_11951_),
    .Y(_11952_));
 sky130_fd_sc_hd__a21oi_1 _18663_ (.A1(_11822_),
    .A2(_11948_),
    .B1(_11952_),
    .Y(_11953_));
 sky130_fd_sc_hd__buf_2 _18664_ (.A(_11699_),
    .X(_11954_));
 sky130_fd_sc_hd__nand2_1 _18665_ (.A(_10626_),
    .B(_11954_),
    .Y(_11955_));
 sky130_fd_sc_hd__xnor2_1 _18666_ (.A(_11953_),
    .B(_11955_),
    .Y(_11956_));
 sky130_fd_sc_hd__clkbuf_2 _18667_ (.A(\genblk1.pcpi_mul.rs1[19] ),
    .X(_11957_));
 sky130_fd_sc_hd__buf_2 _18668_ (.A(_11957_),
    .X(_11958_));
 sky130_fd_sc_hd__buf_2 _18669_ (.A(_11958_),
    .X(_11959_));
 sky130_fd_sc_hd__nand2_1 _18670_ (.A(_10669_),
    .B(_11959_),
    .Y(_11960_));
 sky130_fd_sc_hd__clkbuf_4 _18671_ (.A(_11488_),
    .X(_11961_));
 sky130_fd_sc_hd__and4_1 _18672_ (.A(_11063_),
    .B(_10708_),
    .C(_11380_),
    .D(_11961_),
    .X(_11962_));
 sky130_fd_sc_hd__a22oi_1 _18673_ (.A1(_11058_),
    .A2(_11834_),
    .B1(_11825_),
    .B2(_10662_),
    .Y(_11963_));
 sky130_fd_sc_hd__nor2_1 _18674_ (.A(_11962_),
    .B(_11963_),
    .Y(_11964_));
 sky130_fd_sc_hd__xnor2_2 _18675_ (.A(_11960_),
    .B(_11964_),
    .Y(_11965_));
 sky130_fd_sc_hd__o21ba_1 _18676_ (.A1(_11832_),
    .A2(_11835_),
    .B1_N(_11833_),
    .X(_11966_));
 sky130_fd_sc_hd__xnor2_1 _18677_ (.A(_11965_),
    .B(_11966_),
    .Y(_11967_));
 sky130_fd_sc_hd__xnor2_1 _18678_ (.A(_11956_),
    .B(_11967_),
    .Y(_11968_));
 sky130_fd_sc_hd__a21oi_1 _18679_ (.A1(_11943_),
    .A2(_11944_),
    .B1(_11968_),
    .Y(_11969_));
 sky130_fd_sc_hd__and3_1 _18680_ (.A(_11943_),
    .B(_11944_),
    .C(_11968_),
    .X(_11970_));
 sky130_fd_sc_hd__a211oi_1 _18681_ (.A1(_11941_),
    .A2(_11942_),
    .B1(_11969_),
    .C1(_11970_),
    .Y(_11971_));
 sky130_fd_sc_hd__o211a_1 _18682_ (.A1(_11969_),
    .A2(_11970_),
    .B1(_11941_),
    .C1(_11942_),
    .X(_11972_));
 sky130_fd_sc_hd__nand3_1 _18683_ (.A(_11845_),
    .B(_11855_),
    .C(_11856_),
    .Y(_11973_));
 sky130_fd_sc_hd__a21o_1 _18684_ (.A1(_11793_),
    .A2(_11802_),
    .B1(_11801_),
    .X(_11974_));
 sky130_fd_sc_hd__nand2_1 _18685_ (.A(_11849_),
    .B(_11851_),
    .Y(_11975_));
 sky130_fd_sc_hd__a31o_1 _18686_ (.A1(_10893_),
    .A2(_11037_),
    .A3(_11791_),
    .B1(_11790_),
    .X(_11976_));
 sky130_fd_sc_hd__nand4_2 _18687_ (.A(_11084_),
    .B(_11086_),
    .C(_11067_),
    .D(_11601_),
    .Y(_11977_));
 sky130_fd_sc_hd__a22o_1 _18688_ (.A1(_11196_),
    .A2(_11067_),
    .B1(_11171_),
    .B2(_11298_),
    .X(_11978_));
 sky130_fd_sc_hd__nand4_2 _18689_ (.A(_11089_),
    .B(_11479_),
    .C(_11977_),
    .D(_11978_),
    .Y(_11979_));
 sky130_fd_sc_hd__a22o_1 _18690_ (.A1(_11089_),
    .A2(_11479_),
    .B1(_11977_),
    .B2(_11978_),
    .X(_11980_));
 sky130_fd_sc_hd__nand3_2 _18691_ (.A(_11976_),
    .B(_11979_),
    .C(_11980_),
    .Y(_11981_));
 sky130_fd_sc_hd__a21o_1 _18692_ (.A1(_11979_),
    .A2(_11980_),
    .B1(_11976_),
    .X(_11982_));
 sky130_fd_sc_hd__nand3_2 _18693_ (.A(_11975_),
    .B(_11981_),
    .C(_11982_),
    .Y(_11983_));
 sky130_fd_sc_hd__a21o_1 _18694_ (.A1(_11981_),
    .A2(_11982_),
    .B1(_11975_),
    .X(_11984_));
 sky130_fd_sc_hd__and3_2 _18695_ (.A(_11974_),
    .B(_11983_),
    .C(_11984_),
    .X(_11985_));
 sky130_fd_sc_hd__a21oi_2 _18696_ (.A1(_11983_),
    .A2(_11984_),
    .B1(_11974_),
    .Y(_11986_));
 sky130_fd_sc_hd__a211oi_4 _18697_ (.A1(_11853_),
    .A2(_11855_),
    .B1(_11985_),
    .C1(_11986_),
    .Y(_11987_));
 sky130_fd_sc_hd__o211a_1 _18698_ (.A1(_11985_),
    .A2(_11986_),
    .B1(_11853_),
    .C1(_11855_),
    .X(_11988_));
 sky130_fd_sc_hd__a211oi_2 _18699_ (.A1(_11973_),
    .A2(_11859_),
    .B1(_11987_),
    .C1(_11988_),
    .Y(_11989_));
 sky130_fd_sc_hd__o211a_1 _18700_ (.A1(_11987_),
    .A2(_11988_),
    .B1(_11973_),
    .C1(_11859_),
    .X(_11990_));
 sky130_fd_sc_hd__nor4_1 _18701_ (.A(_11971_),
    .B(_11972_),
    .C(_11989_),
    .D(_11990_),
    .Y(_11991_));
 sky130_fd_sc_hd__o22a_1 _18702_ (.A1(_11971_),
    .A2(_11972_),
    .B1(_11989_),
    .B2(_11990_),
    .X(_11992_));
 sky130_fd_sc_hd__nor3_1 _18703_ (.A(_11807_),
    .B(net357),
    .C(_11992_),
    .Y(_11993_));
 sky130_fd_sc_hd__o21a_1 _18704_ (.A1(net358),
    .A2(_11992_),
    .B1(_11807_),
    .X(_11994_));
 sky130_fd_sc_hd__a211o_1 _18705_ (.A1(_11861_),
    .A2(_11863_),
    .B1(_11993_),
    .C1(_11994_),
    .X(_11995_));
 sky130_fd_sc_hd__o211ai_2 _18706_ (.A1(_11993_),
    .A2(_11994_),
    .B1(_11861_),
    .C1(_11863_),
    .Y(_11996_));
 sky130_fd_sc_hd__nand3_2 _18707_ (.A(_11940_),
    .B(_11995_),
    .C(_11996_),
    .Y(_11997_));
 sky130_fd_sc_hd__a21o_1 _18708_ (.A1(_11995_),
    .A2(_11996_),
    .B1(_11940_),
    .X(_11998_));
 sky130_fd_sc_hd__and3_1 _18709_ (.A(_11869_),
    .B(_11997_),
    .C(_11998_),
    .X(_11999_));
 sky130_fd_sc_hd__a21oi_1 _18710_ (.A1(_11997_),
    .A2(_11998_),
    .B1(_11869_),
    .Y(_12000_));
 sky130_fd_sc_hd__nor3_1 _18711_ (.A(_11888_),
    .B(_11999_),
    .C(_12000_),
    .Y(_12001_));
 sky130_fd_sc_hd__o21a_1 _18712_ (.A1(_11999_),
    .A2(_12000_),
    .B1(_11888_),
    .X(_12002_));
 sky130_fd_sc_hd__a211oi_1 _18713_ (.A1(_11871_),
    .A2(_11885_),
    .B1(net338),
    .C1(_12002_),
    .Y(_12003_));
 sky130_fd_sc_hd__o211a_1 _18714_ (.A1(net338),
    .A2(_12002_),
    .B1(_11871_),
    .C1(_11885_),
    .X(_12004_));
 sky130_fd_sc_hd__or3_2 _18715_ (.A(_11884_),
    .B(_12003_),
    .C(_12004_),
    .X(_12005_));
 sky130_fd_sc_hd__o21ai_1 _18716_ (.A1(_12003_),
    .A2(_12004_),
    .B1(_11884_),
    .Y(_12006_));
 sky130_fd_sc_hd__a211oi_1 _18717_ (.A1(_12005_),
    .A2(_12006_),
    .B1(_11875_),
    .C1(net337),
    .Y(_12007_));
 sky130_fd_sc_hd__o211a_1 _18718_ (.A1(_11875_),
    .A2(net337),
    .B1(_12005_),
    .C1(_12006_),
    .X(_12008_));
 sky130_fd_sc_hd__nor2_1 _18719_ (.A(_12007_),
    .B(_12008_),
    .Y(_12009_));
 sky130_fd_sc_hd__a21oi_1 _18720_ (.A1(_11881_),
    .A2(_11883_),
    .B1(_11879_),
    .Y(_12010_));
 sky130_fd_sc_hd__xnor2_1 _18721_ (.A(_12009_),
    .B(_12010_),
    .Y(_00065_));
 sky130_vsdinv _18722_ (.A(_12003_),
    .Y(_12011_));
 sky130_fd_sc_hd__or2_1 _18723_ (.A(_11886_),
    .B(_11887_),
    .X(_12012_));
 sky130_fd_sc_hd__or3_1 _18724_ (.A(_11807_),
    .B(net357),
    .C(_11992_),
    .X(_12013_));
 sky130_fd_sc_hd__nor2_1 _18725_ (.A(_11969_),
    .B(_11971_),
    .Y(_12014_));
 sky130_fd_sc_hd__a21o_1 _18726_ (.A1(_12013_),
    .A2(_11995_),
    .B1(_12014_),
    .X(_12015_));
 sky130_fd_sc_hd__nand3_1 _18727_ (.A(_12013_),
    .B(_11995_),
    .C(_12014_),
    .Y(_12016_));
 sky130_fd_sc_hd__nand2_1 _18728_ (.A(_12015_),
    .B(_12016_),
    .Y(_12017_));
 sky130_fd_sc_hd__or2_1 _18729_ (.A(_11810_),
    .B(_11939_),
    .X(_12018_));
 sky130_fd_sc_hd__nand2_2 _18730_ (.A(_11778_),
    .B(_11770_),
    .Y(_12019_));
 sky130_fd_sc_hd__clkbuf_2 _18731_ (.A(\genblk1.pcpi_mul.rs2[20] ),
    .X(_12020_));
 sky130_fd_sc_hd__buf_2 _18732_ (.A(_12020_),
    .X(_12021_));
 sky130_fd_sc_hd__and4_1 _18733_ (.A(_10588_),
    .B(_10635_),
    .C(_11890_),
    .D(_12021_),
    .X(_12022_));
 sky130_fd_sc_hd__buf_2 _18734_ (.A(_12021_),
    .X(_12023_));
 sky130_fd_sc_hd__a22oi_2 _18735_ (.A1(_10595_),
    .A2(_11890_),
    .B1(_12023_),
    .B2(_10588_),
    .Y(_12024_));
 sky130_fd_sc_hd__nor2_2 _18736_ (.A(_12022_),
    .B(_12024_),
    .Y(_12025_));
 sky130_fd_sc_hd__xnor2_4 _18737_ (.A(_12019_),
    .B(_12025_),
    .Y(_12026_));
 sky130_fd_sc_hd__nand2_1 _18738_ (.A(_11920_),
    .B(_11932_),
    .Y(_12027_));
 sky130_fd_sc_hd__nand2_1 _18739_ (.A(_11900_),
    .B(_11160_),
    .Y(_12028_));
 sky130_fd_sc_hd__and4_1 _18740_ (.A(_10968_),
    .B(_10962_),
    .C(_11154_),
    .D(_11110_),
    .X(_12029_));
 sky130_fd_sc_hd__a22o_1 _18741_ (.A1(_11904_),
    .A2(_10976_),
    .B1(_11905_),
    .B2(_10968_),
    .X(_12030_));
 sky130_fd_sc_hd__and2b_1 _18742_ (.A_N(_12029_),
    .B(_12030_),
    .X(_12031_));
 sky130_fd_sc_hd__xnor2_1 _18743_ (.A(_12028_),
    .B(_12031_),
    .Y(_12032_));
 sky130_fd_sc_hd__nand2_1 _18744_ (.A(_10858_),
    .B(_11134_),
    .Y(_12033_));
 sky130_fd_sc_hd__and4_1 _18745_ (.A(_10978_),
    .B(_10849_),
    .C(_11240_),
    .D(_11910_),
    .X(_12034_));
 sky130_fd_sc_hd__a22oi_2 _18746_ (.A1(_10909_),
    .A2(_11795_),
    .B1(_11455_),
    .B2(_10848_),
    .Y(_12035_));
 sky130_fd_sc_hd__or3_1 _18747_ (.A(_12033_),
    .B(_12034_),
    .C(_12035_),
    .X(_12036_));
 sky130_fd_sc_hd__o21ai_1 _18748_ (.A1(_12034_),
    .A2(_12035_),
    .B1(_12033_),
    .Y(_12037_));
 sky130_fd_sc_hd__o21bai_1 _18749_ (.A1(_11909_),
    .A2(_11912_),
    .B1_N(_11911_),
    .Y(_12038_));
 sky130_fd_sc_hd__and3_1 _18750_ (.A(_12036_),
    .B(_12037_),
    .C(_12038_),
    .X(_12039_));
 sky130_fd_sc_hd__a21o_1 _18751_ (.A1(_12036_),
    .A2(_12037_),
    .B1(_12038_),
    .X(_12040_));
 sky130_fd_sc_hd__and2b_1 _18752_ (.A_N(_12039_),
    .B(_12040_),
    .X(_12041_));
 sky130_fd_sc_hd__xnor2_1 _18753_ (.A(_12032_),
    .B(_12041_),
    .Y(_12042_));
 sky130_fd_sc_hd__and2b_1 _18754_ (.A_N(_11931_),
    .B(_11930_),
    .X(_12043_));
 sky130_fd_sc_hd__a31o_2 _18755_ (.A1(_10667_),
    .A2(_11445_),
    .A3(_11929_),
    .B1(_11926_),
    .X(_12044_));
 sky130_fd_sc_hd__nand2_1 _18756_ (.A(_11199_),
    .B(_11559_),
    .Y(_12045_));
 sky130_fd_sc_hd__and4_1 _18757_ (.A(_10717_),
    .B(_10719_),
    .C(_11922_),
    .D(_11924_),
    .X(_12046_));
 sky130_fd_sc_hd__a22oi_1 _18758_ (.A1(_10744_),
    .A2(_11555_),
    .B1(_11781_),
    .B2(_10675_),
    .Y(_12047_));
 sky130_fd_sc_hd__nor2_1 _18759_ (.A(_12046_),
    .B(_12047_),
    .Y(_12048_));
 sky130_fd_sc_hd__xnor2_2 _18760_ (.A(_12045_),
    .B(_12048_),
    .Y(_12049_));
 sky130_fd_sc_hd__xnor2_1 _18761_ (.A(_11897_),
    .B(_12049_),
    .Y(_12050_));
 sky130_fd_sc_hd__xnor2_1 _18762_ (.A(_12044_),
    .B(_12050_),
    .Y(_12051_));
 sky130_fd_sc_hd__xnor2_1 _18763_ (.A(_12043_),
    .B(_12051_),
    .Y(_12052_));
 sky130_fd_sc_hd__nor2_1 _18764_ (.A(_12042_),
    .B(_12052_),
    .Y(_12053_));
 sky130_fd_sc_hd__and2_1 _18765_ (.A(_12042_),
    .B(_12052_),
    .X(_12054_));
 sky130_fd_sc_hd__a211o_1 _18766_ (.A1(_12027_),
    .A2(_11934_),
    .B1(_12053_),
    .C1(_12054_),
    .X(_12055_));
 sky130_fd_sc_hd__o211ai_2 _18767_ (.A1(_12053_),
    .A2(_12054_),
    .B1(_12027_),
    .C1(_11934_),
    .Y(_12056_));
 sky130_fd_sc_hd__and3_1 _18768_ (.A(_12026_),
    .B(_12055_),
    .C(_12056_),
    .X(_12057_));
 sky130_fd_sc_hd__a21oi_1 _18769_ (.A1(_12055_),
    .A2(_12056_),
    .B1(_12026_),
    .Y(_12058_));
 sky130_fd_sc_hd__nand2_1 _18770_ (.A(_11898_),
    .B(_11938_),
    .Y(_12059_));
 sky130_fd_sc_hd__o21a_1 _18771_ (.A1(_12057_),
    .A2(_12058_),
    .B1(_12059_),
    .X(_12060_));
 sky130_fd_sc_hd__nor3_1 _18772_ (.A(_12059_),
    .B(_12057_),
    .C(_12058_),
    .Y(_12061_));
 sky130_fd_sc_hd__nor2_1 _18773_ (.A(_11989_),
    .B(_11991_),
    .Y(_12062_));
 sky130_fd_sc_hd__or2_1 _18774_ (.A(_11821_),
    .B(_11951_),
    .X(_12063_));
 sky130_fd_sc_hd__a211o_1 _18775_ (.A1(_11822_),
    .A2(_11948_),
    .B1(_11955_),
    .C1(_11952_),
    .X(_12064_));
 sky130_fd_sc_hd__or2b_1 _18776_ (.A(_11966_),
    .B_N(_11965_),
    .X(_12065_));
 sky130_fd_sc_hd__nand2_1 _18777_ (.A(_11956_),
    .B(_11967_),
    .Y(_12066_));
 sky130_fd_sc_hd__clkbuf_4 _18778_ (.A(_11957_),
    .X(_12067_));
 sky130_fd_sc_hd__nand2_2 _18779_ (.A(_10640_),
    .B(_12067_),
    .Y(_12068_));
 sky130_fd_sc_hd__clkbuf_2 _18780_ (.A(\genblk1.pcpi_mul.rs1[19] ),
    .X(_12069_));
 sky130_fd_sc_hd__clkbuf_4 _18781_ (.A(_12069_),
    .X(_12070_));
 sky130_fd_sc_hd__nand2_1 _18782_ (.A(_10611_),
    .B(_12070_),
    .Y(_12071_));
 sky130_fd_sc_hd__nor2_1 _18783_ (.A(_11948_),
    .B(_12071_),
    .Y(_12072_));
 sky130_fd_sc_hd__a21oi_1 _18784_ (.A1(_11951_),
    .A2(_12068_),
    .B1(_12072_),
    .Y(_12073_));
 sky130_fd_sc_hd__clkbuf_4 _18785_ (.A(_11818_),
    .X(_12074_));
 sky130_fd_sc_hd__buf_4 _18786_ (.A(_12074_),
    .X(_12075_));
 sky130_fd_sc_hd__nand2_2 _18787_ (.A(_11704_),
    .B(_12075_),
    .Y(_12076_));
 sky130_fd_sc_hd__xnor2_1 _18788_ (.A(_12073_),
    .B(_12076_),
    .Y(_12077_));
 sky130_fd_sc_hd__buf_2 _18789_ (.A(\genblk1.pcpi_mul.rs1[20] ),
    .X(_12078_));
 sky130_fd_sc_hd__clkbuf_4 _18790_ (.A(_12078_),
    .X(_12079_));
 sky130_fd_sc_hd__nand2_1 _18791_ (.A(_10669_),
    .B(_12079_),
    .Y(_12080_));
 sky130_fd_sc_hd__clkbuf_2 _18792_ (.A(_11697_),
    .X(_12081_));
 sky130_fd_sc_hd__and4_1 _18793_ (.A(_11710_),
    .B(_10702_),
    .C(_11589_),
    .D(_12081_),
    .X(_12082_));
 sky130_fd_sc_hd__a22oi_1 _18794_ (.A1(_10708_),
    .A2(_11489_),
    .B1(_11598_),
    .B2(_11063_),
    .Y(_12083_));
 sky130_fd_sc_hd__nor2_1 _18795_ (.A(_12082_),
    .B(_12083_),
    .Y(_12084_));
 sky130_fd_sc_hd__xnor2_2 _18796_ (.A(_12080_),
    .B(_12084_),
    .Y(_12085_));
 sky130_fd_sc_hd__o21ba_2 _18797_ (.A1(_11960_),
    .A2(_11963_),
    .B1_N(_11962_),
    .X(_12086_));
 sky130_fd_sc_hd__xnor2_1 _18798_ (.A(_12085_),
    .B(_12086_),
    .Y(_12087_));
 sky130_fd_sc_hd__xnor2_1 _18799_ (.A(_12077_),
    .B(_12087_),
    .Y(_12088_));
 sky130_fd_sc_hd__a21oi_1 _18800_ (.A1(_12065_),
    .A2(_12066_),
    .B1(_12088_),
    .Y(_12089_));
 sky130_fd_sc_hd__and3_1 _18801_ (.A(_12065_),
    .B(_12066_),
    .C(_12088_),
    .X(_12090_));
 sky130_fd_sc_hd__a211oi_1 _18802_ (.A1(_12063_),
    .A2(_12064_),
    .B1(_12089_),
    .C1(_12090_),
    .Y(_12091_));
 sky130_fd_sc_hd__o211a_1 _18803_ (.A1(_12089_),
    .A2(_12090_),
    .B1(_12063_),
    .C1(_12064_),
    .X(_12092_));
 sky130_fd_sc_hd__a21o_1 _18804_ (.A1(_11908_),
    .A2(_11917_),
    .B1(_11916_),
    .X(_12093_));
 sky130_fd_sc_hd__nand2_2 _18805_ (.A(_11977_),
    .B(_11979_),
    .Y(_12094_));
 sky130_fd_sc_hd__a31o_1 _18806_ (.A1(_10892_),
    .A2(_11269_),
    .A3(_11906_),
    .B1(_11902_),
    .X(_12095_));
 sky130_fd_sc_hd__nand2_1 _18807_ (.A(_10787_),
    .B(_11476_),
    .Y(_12096_));
 sky130_fd_sc_hd__nand4_2 _18808_ (.A(_10782_),
    .B(_11200_),
    .C(_11260_),
    .D(_11276_),
    .Y(_12097_));
 sky130_fd_sc_hd__buf_2 _18809_ (.A(\genblk1.pcpi_mul.rs1[12] ),
    .X(_12098_));
 sky130_fd_sc_hd__a22o_1 _18810_ (.A1(_11085_),
    .A2(_12098_),
    .B1(_11371_),
    .B2(_10997_),
    .X(_12099_));
 sky130_fd_sc_hd__nand3b_1 _18811_ (.A_N(_12096_),
    .B(_12097_),
    .C(_12099_),
    .Y(_12100_));
 sky130_fd_sc_hd__a21bo_1 _18812_ (.A1(_12097_),
    .A2(_12099_),
    .B1_N(_12096_),
    .X(_12101_));
 sky130_fd_sc_hd__nand3_2 _18813_ (.A(_12095_),
    .B(_12100_),
    .C(_12101_),
    .Y(_12102_));
 sky130_fd_sc_hd__a21o_1 _18814_ (.A1(_12100_),
    .A2(_12101_),
    .B1(_12095_),
    .X(_12103_));
 sky130_fd_sc_hd__nand3_2 _18815_ (.A(_12094_),
    .B(_12102_),
    .C(_12103_),
    .Y(_12104_));
 sky130_fd_sc_hd__a21o_1 _18816_ (.A1(_12102_),
    .A2(_12103_),
    .B1(_12094_),
    .X(_12105_));
 sky130_fd_sc_hd__and3_1 _18817_ (.A(_12093_),
    .B(_12104_),
    .C(_12105_),
    .X(_12106_));
 sky130_fd_sc_hd__a21oi_2 _18818_ (.A1(_12104_),
    .A2(_12105_),
    .B1(_12093_),
    .Y(_12107_));
 sky130_fd_sc_hd__a211o_2 _18819_ (.A1(_11981_),
    .A2(_11983_),
    .B1(_12106_),
    .C1(_12107_),
    .X(_12108_));
 sky130_fd_sc_hd__o211ai_2 _18820_ (.A1(_12106_),
    .A2(_12107_),
    .B1(_11981_),
    .C1(_11983_),
    .Y(_12109_));
 sky130_fd_sc_hd__o211ai_4 _18821_ (.A1(_11985_),
    .A2(_11987_),
    .B1(_12108_),
    .C1(_12109_),
    .Y(_12110_));
 sky130_fd_sc_hd__a211o_1 _18822_ (.A1(_12108_),
    .A2(_12109_),
    .B1(_11985_),
    .C1(_11987_),
    .X(_12111_));
 sky130_fd_sc_hd__or4bb_2 _18823_ (.A(_12091_),
    .B(_12092_),
    .C_N(_12110_),
    .D_N(_12111_),
    .X(_12112_));
 sky130_fd_sc_hd__a2bb2o_1 _18824_ (.A1_N(_12091_),
    .A2_N(_12092_),
    .B1(_12110_),
    .B2(_12111_),
    .X(_12113_));
 sky130_fd_sc_hd__and3_1 _18825_ (.A(_11936_),
    .B(_12112_),
    .C(_12113_),
    .X(_12114_));
 sky130_fd_sc_hd__a21oi_1 _18826_ (.A1(_12112_),
    .A2(_12113_),
    .B1(_11936_),
    .Y(_12115_));
 sky130_fd_sc_hd__nor3_1 _18827_ (.A(_12062_),
    .B(_12114_),
    .C(_12115_),
    .Y(_12116_));
 sky130_fd_sc_hd__o21a_1 _18828_ (.A1(_12114_),
    .A2(_12115_),
    .B1(_12062_),
    .X(_12117_));
 sky130_fd_sc_hd__nor4_2 _18829_ (.A(_12060_),
    .B(net343),
    .C(_12116_),
    .D(_12117_),
    .Y(_12118_));
 sky130_fd_sc_hd__o22a_1 _18830_ (.A1(_12060_),
    .A2(net343),
    .B1(_12116_),
    .B2(_12117_),
    .X(_12119_));
 sky130_fd_sc_hd__a211oi_2 _18831_ (.A1(_12018_),
    .A2(_11997_),
    .B1(net339),
    .C1(_12119_),
    .Y(_12120_));
 sky130_fd_sc_hd__o211a_1 _18832_ (.A1(net339),
    .A2(_12119_),
    .B1(_12018_),
    .C1(_11997_),
    .X(_12121_));
 sky130_fd_sc_hd__or3_1 _18833_ (.A(_12017_),
    .B(_12120_),
    .C(_12121_),
    .X(_12122_));
 sky130_fd_sc_hd__o21ai_1 _18834_ (.A1(_12120_),
    .A2(_12121_),
    .B1(_12017_),
    .Y(_12123_));
 sky130_fd_sc_hd__o211a_1 _18835_ (.A1(_11999_),
    .A2(_12001_),
    .B1(_12122_),
    .C1(_12123_),
    .X(_12124_));
 sky130_fd_sc_hd__a211oi_1 _18836_ (.A1(_12122_),
    .A2(_12123_),
    .B1(_11999_),
    .C1(_12001_),
    .Y(_12125_));
 sky130_fd_sc_hd__nor3_1 _18837_ (.A(_12012_),
    .B(_12124_),
    .C(_12125_),
    .Y(_12126_));
 sky130_fd_sc_hd__o21a_1 _18838_ (.A1(_12124_),
    .A2(_12125_),
    .B1(_12012_),
    .X(_12127_));
 sky130_fd_sc_hd__a211oi_1 _18839_ (.A1(_12011_),
    .A2(_12005_),
    .B1(_12126_),
    .C1(_12127_),
    .Y(_12128_));
 sky130_fd_sc_hd__o211a_1 _18840_ (.A1(_12126_),
    .A2(_12127_),
    .B1(_12011_),
    .C1(_12005_),
    .X(_12129_));
 sky130_fd_sc_hd__or2_1 _18841_ (.A(_12128_),
    .B(_12129_),
    .X(_12130_));
 sky130_fd_sc_hd__nand4b_1 _18842_ (.A_N(_11645_),
    .B(_11761_),
    .C(_11881_),
    .D(_12009_),
    .Y(_12131_));
 sky130_fd_sc_hd__and2b_1 _18843_ (.A_N(_12007_),
    .B(_11879_),
    .X(_12132_));
 sky130_fd_sc_hd__a311o_1 _18844_ (.A1(_11881_),
    .A2(_11882_),
    .A3(_12009_),
    .B1(_12132_),
    .C1(_12008_),
    .X(_12133_));
 sky130_fd_sc_hd__o21ba_1 _18845_ (.A1(_11548_),
    .A2(_12131_),
    .B1_N(_12133_),
    .X(_12134_));
 sky130_fd_sc_hd__xor2_1 _18846_ (.A(_12130_),
    .B(_12134_),
    .X(_00066_));
 sky130_fd_sc_hd__nor3_1 _18847_ (.A(_12017_),
    .B(_12120_),
    .C(_12121_),
    .Y(_12135_));
 sky130_fd_sc_hd__nor2_1 _18848_ (.A(_12114_),
    .B(_12116_),
    .Y(_12136_));
 sky130_fd_sc_hd__nor2_1 _18849_ (.A(_12089_),
    .B(_12091_),
    .Y(_12137_));
 sky130_fd_sc_hd__xnor2_1 _18850_ (.A(_12136_),
    .B(_12137_),
    .Y(_12138_));
 sky130_fd_sc_hd__or2_1 _18851_ (.A(_11948_),
    .B(_12071_),
    .X(_12139_));
 sky130_fd_sc_hd__a211o_1 _18852_ (.A1(_11951_),
    .A2(_12068_),
    .B1(_12076_),
    .C1(_12072_),
    .X(_12140_));
 sky130_fd_sc_hd__or2b_1 _18853_ (.A(_12086_),
    .B_N(_12085_),
    .X(_12141_));
 sky130_fd_sc_hd__nand2_1 _18854_ (.A(_12077_),
    .B(_12087_),
    .Y(_12142_));
 sky130_fd_sc_hd__clkbuf_2 _18855_ (.A(\genblk1.pcpi_mul.rs1[20] ),
    .X(_12143_));
 sky130_fd_sc_hd__buf_2 _18856_ (.A(_12143_),
    .X(_12144_));
 sky130_fd_sc_hd__clkbuf_4 _18857_ (.A(_12144_),
    .X(_12145_));
 sky130_fd_sc_hd__nand2_4 _18858_ (.A(_10600_),
    .B(_12145_),
    .Y(_12146_));
 sky130_fd_sc_hd__buf_4 _18859_ (.A(_12078_),
    .X(_12147_));
 sky130_fd_sc_hd__nand2_1 _18860_ (.A(_10740_),
    .B(_12147_),
    .Y(_12148_));
 sky130_fd_sc_hd__nor2_1 _18861_ (.A(_12068_),
    .B(_12148_),
    .Y(_12149_));
 sky130_fd_sc_hd__a21oi_1 _18862_ (.A1(_12071_),
    .A2(_12146_),
    .B1(_12149_),
    .Y(_12150_));
 sky130_fd_sc_hd__nand2_2 _18863_ (.A(_10625_),
    .B(_11950_),
    .Y(_12151_));
 sky130_fd_sc_hd__xnor2_1 _18864_ (.A(_12150_),
    .B(_12151_),
    .Y(_12152_));
 sky130_fd_sc_hd__clkbuf_2 _18865_ (.A(\genblk1.pcpi_mul.rs1[21] ),
    .X(_12153_));
 sky130_fd_sc_hd__clkbuf_4 _18866_ (.A(_12153_),
    .X(_12154_));
 sky130_fd_sc_hd__nand2_1 _18867_ (.A(_10583_),
    .B(_12154_),
    .Y(_12155_));
 sky130_fd_sc_hd__and4_1 _18868_ (.A(_10661_),
    .B(_10707_),
    .C(_11597_),
    .D(_11818_),
    .X(_12156_));
 sky130_fd_sc_hd__a22oi_2 _18869_ (.A1(_10702_),
    .A2(_12081_),
    .B1(_11707_),
    .B2(_11710_),
    .Y(_12157_));
 sky130_fd_sc_hd__nor2_1 _18870_ (.A(_12156_),
    .B(_12157_),
    .Y(_12158_));
 sky130_fd_sc_hd__xnor2_2 _18871_ (.A(_12155_),
    .B(_12158_),
    .Y(_12159_));
 sky130_fd_sc_hd__o21ba_1 _18872_ (.A1(_12080_),
    .A2(_12083_),
    .B1_N(_12082_),
    .X(_12160_));
 sky130_fd_sc_hd__xnor2_1 _18873_ (.A(_12159_),
    .B(_12160_),
    .Y(_12161_));
 sky130_fd_sc_hd__xnor2_1 _18874_ (.A(_12152_),
    .B(_12161_),
    .Y(_12162_));
 sky130_fd_sc_hd__a21oi_1 _18875_ (.A1(_12141_),
    .A2(_12142_),
    .B1(_12162_),
    .Y(_12163_));
 sky130_fd_sc_hd__and3_1 _18876_ (.A(_12141_),
    .B(_12142_),
    .C(_12162_),
    .X(_12164_));
 sky130_fd_sc_hd__a211oi_1 _18877_ (.A1(_12139_),
    .A2(_12140_),
    .B1(_12163_),
    .C1(_12164_),
    .Y(_12165_));
 sky130_fd_sc_hd__o211a_1 _18878_ (.A1(_12163_),
    .A2(_12164_),
    .B1(_12139_),
    .C1(_12140_),
    .X(_12166_));
 sky130_fd_sc_hd__nand3_1 _18879_ (.A(_12093_),
    .B(_12104_),
    .C(_12105_),
    .Y(_12167_));
 sky130_fd_sc_hd__a21o_1 _18880_ (.A1(_12032_),
    .A2(_12040_),
    .B1(_12039_),
    .X(_12168_));
 sky130_fd_sc_hd__nand2_1 _18881_ (.A(_12097_),
    .B(_12100_),
    .Y(_12169_));
 sky130_fd_sc_hd__a31o_1 _18882_ (.A1(_10960_),
    .A2(_11055_),
    .A3(_12030_),
    .B1(_12029_),
    .X(_12170_));
 sky130_fd_sc_hd__nand4_2 _18883_ (.A(_10782_),
    .B(_11200_),
    .C(_11276_),
    .D(_11481_),
    .Y(_12171_));
 sky130_fd_sc_hd__buf_2 _18884_ (.A(_10781_),
    .X(_12172_));
 sky130_fd_sc_hd__a22o_1 _18885_ (.A1(_11085_),
    .A2(_11371_),
    .B1(_11379_),
    .B2(_12172_),
    .X(_12173_));
 sky130_fd_sc_hd__nand4_2 _18886_ (.A(_11508_),
    .B(_11590_),
    .C(_12171_),
    .D(_12173_),
    .Y(_12174_));
 sky130_fd_sc_hd__a22o_1 _18887_ (.A1(_10736_),
    .A2(_11961_),
    .B1(_12171_),
    .B2(_12173_),
    .X(_12175_));
 sky130_fd_sc_hd__nand3_2 _18888_ (.A(_12170_),
    .B(_12174_),
    .C(_12175_),
    .Y(_12176_));
 sky130_fd_sc_hd__a21o_1 _18889_ (.A1(_12174_),
    .A2(_12175_),
    .B1(_12170_),
    .X(_12177_));
 sky130_fd_sc_hd__nand3_2 _18890_ (.A(_12169_),
    .B(_12176_),
    .C(_12177_),
    .Y(_12178_));
 sky130_fd_sc_hd__a21o_1 _18891_ (.A1(_12176_),
    .A2(_12177_),
    .B1(_12169_),
    .X(_12179_));
 sky130_fd_sc_hd__and3_1 _18892_ (.A(_12168_),
    .B(_12178_),
    .C(_12179_),
    .X(_12180_));
 sky130_fd_sc_hd__a21oi_1 _18893_ (.A1(_12178_),
    .A2(_12179_),
    .B1(_12168_),
    .Y(_12181_));
 sky130_fd_sc_hd__a211oi_2 _18894_ (.A1(_12102_),
    .A2(_12104_),
    .B1(_12180_),
    .C1(_12181_),
    .Y(_12182_));
 sky130_fd_sc_hd__o211a_1 _18895_ (.A1(_12180_),
    .A2(_12181_),
    .B1(_12102_),
    .C1(_12104_),
    .X(_12183_));
 sky130_fd_sc_hd__a211oi_1 _18896_ (.A1(_12167_),
    .A2(_12108_),
    .B1(_12182_),
    .C1(_12183_),
    .Y(_12184_));
 sky130_fd_sc_hd__o211a_1 _18897_ (.A1(_12182_),
    .A2(_12183_),
    .B1(_12167_),
    .C1(_12108_),
    .X(_12185_));
 sky130_fd_sc_hd__or4_1 _18898_ (.A(_12165_),
    .B(_12166_),
    .C(_12184_),
    .D(_12185_),
    .X(_12186_));
 sky130_fd_sc_hd__o22ai_1 _18899_ (.A1(_12165_),
    .A2(_12166_),
    .B1(_12184_),
    .B2(_12185_),
    .Y(_12187_));
 sky130_fd_sc_hd__and3b_1 _18900_ (.A_N(_12055_),
    .B(_12186_),
    .C(_12187_),
    .X(_12188_));
 sky130_fd_sc_hd__a21boi_1 _18901_ (.A1(_12186_),
    .A2(_12187_),
    .B1_N(_12055_),
    .Y(_12189_));
 sky130_fd_sc_hd__a211oi_1 _18902_ (.A1(_12110_),
    .A2(_12112_),
    .B1(_12188_),
    .C1(_12189_),
    .Y(_12190_));
 sky130_fd_sc_hd__o211a_1 _18903_ (.A1(_12188_),
    .A2(_12189_),
    .B1(_12110_),
    .C1(_12112_),
    .X(_12191_));
 sky130_fd_sc_hd__nand3_1 _18904_ (.A(_12026_),
    .B(_12055_),
    .C(_12056_),
    .Y(_12192_));
 sky130_fd_sc_hd__and2_1 _18905_ (.A(_12043_),
    .B(_12051_),
    .X(_12193_));
 sky130_fd_sc_hd__nand2_1 _18906_ (.A(_11190_),
    .B(_11265_),
    .Y(_12194_));
 sky130_fd_sc_hd__and4_1 _18907_ (.A(_11904_),
    .B(_10976_),
    .C(_11905_),
    .D(_11054_),
    .X(_12195_));
 sky130_fd_sc_hd__a22o_1 _18908_ (.A1(_10976_),
    .A2(_11905_),
    .B1(_11054_),
    .B2(_11904_),
    .X(_12196_));
 sky130_fd_sc_hd__and2b_1 _18909_ (.A_N(_12195_),
    .B(_12196_),
    .X(_12197_));
 sky130_fd_sc_hd__xnor2_1 _18910_ (.A(_12194_),
    .B(_12197_),
    .Y(_12198_));
 sky130_fd_sc_hd__nand2_1 _18911_ (.A(_10919_),
    .B(_11134_),
    .Y(_12199_));
 sky130_fd_sc_hd__and4_1 _18912_ (.A(_10849_),
    .B(_11047_),
    .C(_11795_),
    .D(_11353_),
    .X(_12200_));
 sky130_fd_sc_hd__a22oi_2 _18913_ (.A1(_11174_),
    .A2(_11235_),
    .B1(_11458_),
    .B2(_10909_),
    .Y(_12201_));
 sky130_fd_sc_hd__or3_1 _18914_ (.A(_12199_),
    .B(_12200_),
    .C(_12201_),
    .X(_12202_));
 sky130_fd_sc_hd__o21ai_1 _18915_ (.A1(_12200_),
    .A2(_12201_),
    .B1(_12199_),
    .Y(_12203_));
 sky130_fd_sc_hd__o21bai_1 _18916_ (.A1(_12033_),
    .A2(_12035_),
    .B1_N(_12034_),
    .Y(_12204_));
 sky130_fd_sc_hd__and3_1 _18917_ (.A(_12202_),
    .B(_12203_),
    .C(_12204_),
    .X(_12205_));
 sky130_fd_sc_hd__a21o_1 _18918_ (.A1(_12202_),
    .A2(_12203_),
    .B1(_12204_),
    .X(_12206_));
 sky130_fd_sc_hd__and2b_1 _18919_ (.A_N(_12205_),
    .B(_12206_),
    .X(_12207_));
 sky130_fd_sc_hd__xnor2_1 _18920_ (.A(_12198_),
    .B(_12207_),
    .Y(_12208_));
 sky130_fd_sc_hd__and2_1 _18921_ (.A(_11897_),
    .B(_12049_),
    .X(_12209_));
 sky130_fd_sc_hd__and2b_1 _18922_ (.A_N(_12050_),
    .B(_12044_),
    .X(_12210_));
 sky130_fd_sc_hd__o21ba_1 _18923_ (.A1(_12045_),
    .A2(_12047_),
    .B1_N(_12046_),
    .X(_12211_));
 sky130_fd_sc_hd__o21ba_1 _18924_ (.A1(_12019_),
    .A2(_12024_),
    .B1_N(_12022_),
    .X(_12212_));
 sky130_fd_sc_hd__nand2_1 _18925_ (.A(_11302_),
    .B(_11559_),
    .Y(_12213_));
 sky130_fd_sc_hd__and4_1 _18926_ (.A(_10719_),
    .B(_10794_),
    .C(_11662_),
    .D(_11658_),
    .X(_12214_));
 sky130_fd_sc_hd__a22oi_2 _18927_ (.A1(_10697_),
    .A2(_11555_),
    .B1(_11925_),
    .B2(_10742_),
    .Y(_12215_));
 sky130_fd_sc_hd__nor2_1 _18928_ (.A(_12214_),
    .B(_12215_),
    .Y(_12216_));
 sky130_fd_sc_hd__xnor2_2 _18929_ (.A(_12213_),
    .B(_12216_),
    .Y(_12217_));
 sky130_fd_sc_hd__xnor2_1 _18930_ (.A(_12212_),
    .B(_12217_),
    .Y(_12218_));
 sky130_fd_sc_hd__xnor2_1 _18931_ (.A(_12211_),
    .B(_12218_),
    .Y(_12219_));
 sky130_fd_sc_hd__o21a_1 _18932_ (.A1(_12209_),
    .A2(_12210_),
    .B1(_12219_),
    .X(_12220_));
 sky130_fd_sc_hd__nor3_1 _18933_ (.A(_12209_),
    .B(_12210_),
    .C(_12219_),
    .Y(_12221_));
 sky130_fd_sc_hd__or3_1 _18934_ (.A(_12208_),
    .B(_12220_),
    .C(_12221_),
    .X(_12222_));
 sky130_fd_sc_hd__o21ai_1 _18935_ (.A1(_12220_),
    .A2(_12221_),
    .B1(_12208_),
    .Y(_12223_));
 sky130_fd_sc_hd__o211a_1 _18936_ (.A1(_12193_),
    .A2(_12053_),
    .B1(_12222_),
    .C1(_12223_),
    .X(_12224_));
 sky130_fd_sc_hd__a211oi_1 _18937_ (.A1(_12222_),
    .A2(_12223_),
    .B1(_12193_),
    .C1(_12053_),
    .Y(_12225_));
 sky130_fd_sc_hd__buf_2 _18938_ (.A(\genblk1.pcpi_mul.rs2[21] ),
    .X(_12226_));
 sky130_fd_sc_hd__buf_2 _18939_ (.A(_12226_),
    .X(_12227_));
 sky130_fd_sc_hd__clkbuf_4 _18940_ (.A(_12227_),
    .X(_12228_));
 sky130_fd_sc_hd__clkbuf_4 _18941_ (.A(_12228_),
    .X(_12229_));
 sky130_fd_sc_hd__nand2_1 _18942_ (.A(_10590_),
    .B(_12229_),
    .Y(_12230_));
 sky130_fd_sc_hd__nand2_2 _18943_ (.A(_10649_),
    .B(_11894_),
    .Y(_12231_));
 sky130_fd_sc_hd__clkbuf_2 _18944_ (.A(\genblk1.pcpi_mul.rs2[20] ),
    .X(_12232_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18945_ (.A(_12232_),
    .X(_12233_));
 sky130_fd_sc_hd__and4_1 _18946_ (.A(_10594_),
    .B(_10628_),
    .C(_11889_),
    .D(_12233_),
    .X(_12234_));
 sky130_fd_sc_hd__clkbuf_2 _18947_ (.A(_11889_),
    .X(_12235_));
 sky130_fd_sc_hd__a22oi_2 _18948_ (.A1(_11777_),
    .A2(_12235_),
    .B1(_12021_),
    .B2(_10635_),
    .Y(_12236_));
 sky130_fd_sc_hd__nor2_2 _18949_ (.A(_12234_),
    .B(_12236_),
    .Y(_12237_));
 sky130_fd_sc_hd__xnor2_4 _18950_ (.A(_12231_),
    .B(_12237_),
    .Y(_12238_));
 sky130_fd_sc_hd__xnor2_1 _18951_ (.A(_12230_),
    .B(_12238_),
    .Y(_12239_));
 sky130_fd_sc_hd__nor3b_2 _18952_ (.A(_12224_),
    .B(_12225_),
    .C_N(_12239_),
    .Y(_12240_));
 sky130_fd_sc_hd__o21ba_1 _18953_ (.A1(_12224_),
    .A2(_12225_),
    .B1_N(_12239_),
    .X(_12241_));
 sky130_fd_sc_hd__or3_2 _18954_ (.A(_12192_),
    .B(_12240_),
    .C(_12241_),
    .X(_12242_));
 sky130_fd_sc_hd__o21ai_1 _18955_ (.A1(_12240_),
    .A2(_12241_),
    .B1(_12192_),
    .Y(_12243_));
 sky130_fd_sc_hd__or4bb_4 _18956_ (.A(_12190_),
    .B(_12191_),
    .C_N(_12242_),
    .D_N(_12243_),
    .X(_12244_));
 sky130_fd_sc_hd__a2bb2o_1 _18957_ (.A1_N(_12190_),
    .A2_N(_12191_),
    .B1(_12242_),
    .B2(_12243_),
    .X(_12245_));
 sky130_fd_sc_hd__o211a_1 _18958_ (.A1(_12061_),
    .A2(_12118_),
    .B1(_12244_),
    .C1(_12245_),
    .X(_12246_));
 sky130_fd_sc_hd__a211oi_1 _18959_ (.A1(_12244_),
    .A2(_12245_),
    .B1(_12061_),
    .C1(_12118_),
    .Y(_12247_));
 sky130_fd_sc_hd__or3_1 _18960_ (.A(_12138_),
    .B(_12246_),
    .C(_12247_),
    .X(_12248_));
 sky130_fd_sc_hd__o21ai_1 _18961_ (.A1(_12246_),
    .A2(_12247_),
    .B1(_12138_),
    .Y(_12249_));
 sky130_fd_sc_hd__o211a_1 _18962_ (.A1(_12120_),
    .A2(_12135_),
    .B1(_12248_),
    .C1(_12249_),
    .X(_12250_));
 sky130_fd_sc_hd__a211oi_1 _18963_ (.A1(_12248_),
    .A2(_12249_),
    .B1(_12120_),
    .C1(_12135_),
    .Y(_12251_));
 sky130_fd_sc_hd__or3_1 _18964_ (.A(_12015_),
    .B(_12250_),
    .C(_12251_),
    .X(_12252_));
 sky130_fd_sc_hd__o21ai_1 _18965_ (.A1(_12250_),
    .A2(_12251_),
    .B1(_12015_),
    .Y(_12253_));
 sky130_fd_sc_hd__o211a_1 _18966_ (.A1(_12124_),
    .A2(net336),
    .B1(_12252_),
    .C1(_12253_),
    .X(_12254_));
 sky130_fd_sc_hd__a211oi_1 _18967_ (.A1(_12252_),
    .A2(_12253_),
    .B1(_12124_),
    .C1(net336),
    .Y(_12255_));
 sky130_fd_sc_hd__nor2_1 _18968_ (.A(_12254_),
    .B(_12255_),
    .Y(_12256_));
 sky130_fd_sc_hd__nor2_1 _18969_ (.A(_12130_),
    .B(_12134_),
    .Y(_12257_));
 sky130_fd_sc_hd__nor2_1 _18970_ (.A(_12128_),
    .B(_12257_),
    .Y(_12258_));
 sky130_fd_sc_hd__xnor2_1 _18971_ (.A(_12256_),
    .B(_12258_),
    .Y(_00067_));
 sky130_fd_sc_hd__o21ba_1 _18972_ (.A1(_12128_),
    .A2(_12254_),
    .B1_N(_12255_),
    .X(_12259_));
 sky130_fd_sc_hd__a21oi_1 _18973_ (.A1(_12257_),
    .A2(_12256_),
    .B1(_12259_),
    .Y(_12260_));
 sky130_fd_sc_hd__or2_1 _18974_ (.A(_12136_),
    .B(_12137_),
    .X(_12261_));
 sky130_fd_sc_hd__nor3_1 _18975_ (.A(_12138_),
    .B(_12246_),
    .C(_12247_),
    .Y(_12262_));
 sky130_fd_sc_hd__nor2_1 _18976_ (.A(_12188_),
    .B(_12190_),
    .Y(_12263_));
 sky130_fd_sc_hd__nor2_1 _18977_ (.A(_12163_),
    .B(_12165_),
    .Y(_12264_));
 sky130_fd_sc_hd__xnor2_1 _18978_ (.A(_12263_),
    .B(_12264_),
    .Y(_12265_));
 sky130_fd_sc_hd__and2b_1 _18979_ (.A_N(_12184_),
    .B(_12186_),
    .X(_12266_));
 sky130_fd_sc_hd__or2_1 _18980_ (.A(_12068_),
    .B(_12148_),
    .X(_12267_));
 sky130_fd_sc_hd__a211o_1 _18981_ (.A1(_12071_),
    .A2(_12146_),
    .B1(_12151_),
    .C1(_12149_),
    .X(_12268_));
 sky130_fd_sc_hd__or2b_1 _18982_ (.A(_12160_),
    .B_N(_12159_),
    .X(_12269_));
 sky130_fd_sc_hd__nand2_1 _18983_ (.A(_12152_),
    .B(_12161_),
    .Y(_12270_));
 sky130_fd_sc_hd__buf_4 _18984_ (.A(_12153_),
    .X(_12271_));
 sky130_fd_sc_hd__nand2_1 _18985_ (.A(_10640_),
    .B(_12271_),
    .Y(_12272_));
 sky130_fd_sc_hd__clkbuf_4 _18986_ (.A(\genblk1.pcpi_mul.rs1[21] ),
    .X(_12273_));
 sky130_fd_sc_hd__clkbuf_4 _18987_ (.A(_12273_),
    .X(_12274_));
 sky130_fd_sc_hd__nand2_1 _18988_ (.A(_10611_),
    .B(_12274_),
    .Y(_12275_));
 sky130_fd_sc_hd__nor2_1 _18989_ (.A(_12146_),
    .B(_12275_),
    .Y(_12276_));
 sky130_fd_sc_hd__a21oi_1 _18990_ (.A1(_12148_),
    .A2(_12272_),
    .B1(_12276_),
    .Y(_12277_));
 sky130_fd_sc_hd__buf_2 _18991_ (.A(_12070_),
    .X(_12278_));
 sky130_fd_sc_hd__nand2_2 _18992_ (.A(_11704_),
    .B(_12278_),
    .Y(_12279_));
 sky130_fd_sc_hd__xnor2_1 _18993_ (.A(_12277_),
    .B(_12279_),
    .Y(_12280_));
 sky130_fd_sc_hd__clkbuf_2 _18994_ (.A(\genblk1.pcpi_mul.rs1[22] ),
    .X(_12281_));
 sky130_fd_sc_hd__clkbuf_4 _18995_ (.A(_12281_),
    .X(_12282_));
 sky130_fd_sc_hd__nand2_1 _18996_ (.A(_10669_),
    .B(_12282_),
    .Y(_12283_));
 sky130_fd_sc_hd__and4_1 _18997_ (.A(_11710_),
    .B(_10702_),
    .C(_11818_),
    .D(_11946_),
    .X(_12284_));
 sky130_fd_sc_hd__clkbuf_4 _18998_ (.A(_11818_),
    .X(_12285_));
 sky130_fd_sc_hd__a22oi_2 _18999_ (.A1(_10708_),
    .A2(_12285_),
    .B1(_11949_),
    .B2(_11063_),
    .Y(_12286_));
 sky130_fd_sc_hd__nor2_1 _19000_ (.A(_12284_),
    .B(_12286_),
    .Y(_12287_));
 sky130_fd_sc_hd__xnor2_2 _19001_ (.A(_12283_),
    .B(_12287_),
    .Y(_12288_));
 sky130_fd_sc_hd__o21ba_1 _19002_ (.A1(_12155_),
    .A2(_12157_),
    .B1_N(_12156_),
    .X(_12289_));
 sky130_fd_sc_hd__xnor2_1 _19003_ (.A(_12288_),
    .B(_12289_),
    .Y(_12290_));
 sky130_fd_sc_hd__xnor2_1 _19004_ (.A(_12280_),
    .B(_12290_),
    .Y(_12291_));
 sky130_fd_sc_hd__a21oi_1 _19005_ (.A1(_12269_),
    .A2(_12270_),
    .B1(_12291_),
    .Y(_12292_));
 sky130_fd_sc_hd__and3_1 _19006_ (.A(_12269_),
    .B(_12270_),
    .C(_12291_),
    .X(_12293_));
 sky130_fd_sc_hd__a211oi_1 _19007_ (.A1(_12267_),
    .A2(_12268_),
    .B1(_12292_),
    .C1(_12293_),
    .Y(_12294_));
 sky130_fd_sc_hd__o211a_1 _19008_ (.A1(_12292_),
    .A2(_12293_),
    .B1(_12267_),
    .C1(_12268_),
    .X(_12295_));
 sky130_fd_sc_hd__a21o_1 _19009_ (.A1(_12198_),
    .A2(_12206_),
    .B1(_12205_),
    .X(_12296_));
 sky130_fd_sc_hd__nand2_1 _19010_ (.A(_12171_),
    .B(_12174_),
    .Y(_12297_));
 sky130_fd_sc_hd__a31o_1 _19011_ (.A1(_10892_),
    .A2(_11261_),
    .A3(_12196_),
    .B1(_12195_),
    .X(_12298_));
 sky130_fd_sc_hd__nand2_1 _19012_ (.A(_10787_),
    .B(_11698_),
    .Y(_12299_));
 sky130_fd_sc_hd__nand4_2 _19013_ (.A(_11082_),
    .B(_11200_),
    .C(_11481_),
    .D(_11489_),
    .Y(_12300_));
 sky130_fd_sc_hd__a22o_1 _19014_ (.A1(_11200_),
    .A2(_11481_),
    .B1(_11589_),
    .B2(_10997_),
    .X(_12301_));
 sky130_fd_sc_hd__nand3b_1 _19015_ (.A_N(_12299_),
    .B(_12300_),
    .C(_12301_),
    .Y(_12302_));
 sky130_fd_sc_hd__a21bo_1 _19016_ (.A1(_12300_),
    .A2(_12301_),
    .B1_N(_12299_),
    .X(_12303_));
 sky130_fd_sc_hd__nand3_2 _19017_ (.A(_12298_),
    .B(_12302_),
    .C(_12303_),
    .Y(_12304_));
 sky130_fd_sc_hd__a21o_1 _19018_ (.A1(_12302_),
    .A2(_12303_),
    .B1(_12298_),
    .X(_12305_));
 sky130_fd_sc_hd__nand3_2 _19019_ (.A(_12297_),
    .B(_12304_),
    .C(_12305_),
    .Y(_12306_));
 sky130_fd_sc_hd__a21o_1 _19020_ (.A1(_12304_),
    .A2(_12305_),
    .B1(_12297_),
    .X(_12307_));
 sky130_fd_sc_hd__and3_1 _19021_ (.A(_12296_),
    .B(_12306_),
    .C(_12307_),
    .X(_12308_));
 sky130_fd_sc_hd__a21oi_1 _19022_ (.A1(_12306_),
    .A2(_12307_),
    .B1(_12296_),
    .Y(_12309_));
 sky130_fd_sc_hd__a211o_1 _19023_ (.A1(_12176_),
    .A2(_12178_),
    .B1(_12308_),
    .C1(_12309_),
    .X(_12310_));
 sky130_fd_sc_hd__o211ai_2 _19024_ (.A1(_12308_),
    .A2(_12309_),
    .B1(_12176_),
    .C1(_12178_),
    .Y(_12311_));
 sky130_fd_sc_hd__o211ai_2 _19025_ (.A1(_12180_),
    .A2(_12182_),
    .B1(_12310_),
    .C1(_12311_),
    .Y(_12312_));
 sky130_fd_sc_hd__a211o_1 _19026_ (.A1(_12310_),
    .A2(_12311_),
    .B1(_12180_),
    .C1(_12182_),
    .X(_12313_));
 sky130_fd_sc_hd__or4bb_2 _19027_ (.A(_12294_),
    .B(_12295_),
    .C_N(_12312_),
    .D_N(_12313_),
    .X(_12314_));
 sky130_fd_sc_hd__a2bb2o_1 _19028_ (.A1_N(_12294_),
    .A2_N(_12295_),
    .B1(_12312_),
    .B2(_12313_),
    .X(_12315_));
 sky130_fd_sc_hd__and3_1 _19029_ (.A(_12224_),
    .B(_12314_),
    .C(_12315_),
    .X(_12316_));
 sky130_fd_sc_hd__a21oi_1 _19030_ (.A1(_12314_),
    .A2(_12315_),
    .B1(_12224_),
    .Y(_12317_));
 sky130_fd_sc_hd__nor3_1 _19031_ (.A(_12266_),
    .B(_12316_),
    .C(_12317_),
    .Y(_12318_));
 sky130_fd_sc_hd__o21a_1 _19032_ (.A1(_12316_),
    .A2(_12317_),
    .B1(_12266_),
    .X(_12319_));
 sky130_fd_sc_hd__or2b_1 _19033_ (.A(_12230_),
    .B_N(_12238_),
    .X(_12320_));
 sky130_fd_sc_hd__buf_1 _19034_ (.A(\genblk1.pcpi_mul.rs2[22] ),
    .X(_12321_));
 sky130_fd_sc_hd__buf_2 _19035_ (.A(_12321_),
    .X(_12322_));
 sky130_fd_sc_hd__clkbuf_2 _19036_ (.A(_12322_),
    .X(_12323_));
 sky130_fd_sc_hd__clkbuf_4 _19037_ (.A(_12323_),
    .X(_12324_));
 sky130_fd_sc_hd__buf_4 _19038_ (.A(_12324_),
    .X(_12325_));
 sky130_fd_sc_hd__a22oi_4 _19039_ (.A1(_10596_),
    .A2(_12228_),
    .B1(_12325_),
    .B2(_10590_),
    .Y(_12326_));
 sky130_fd_sc_hd__clkbuf_2 _19040_ (.A(\genblk1.pcpi_mul.rs2[22] ),
    .X(_12327_));
 sky130_fd_sc_hd__clkbuf_2 _19041_ (.A(_12327_),
    .X(_12328_));
 sky130_fd_sc_hd__clkbuf_4 _19042_ (.A(_12328_),
    .X(_12329_));
 sky130_fd_sc_hd__and4_2 _19043_ (.A(_10588_),
    .B(_10595_),
    .C(_12226_),
    .D(_12329_),
    .X(_12330_));
 sky130_fd_sc_hd__nor2_1 _19044_ (.A(_12326_),
    .B(_12330_),
    .Y(_12331_));
 sky130_fd_sc_hd__nand2_2 _19045_ (.A(_10667_),
    .B(_11772_),
    .Y(_12332_));
 sky130_fd_sc_hd__buf_1 _19046_ (.A(\genblk1.pcpi_mul.rs2[19] ),
    .X(_12333_));
 sky130_fd_sc_hd__and4_1 _19047_ (.A(_10606_),
    .B(_10647_),
    .C(_12333_),
    .D(_12232_),
    .X(_12334_));
 sky130_fd_sc_hd__a22o_1 _19048_ (.A1(_10800_),
    .A2(_12333_),
    .B1(_12020_),
    .B2(_10606_),
    .X(_12335_));
 sky130_fd_sc_hd__and2b_1 _19049_ (.A_N(_12334_),
    .B(_12335_),
    .X(_12336_));
 sky130_fd_sc_hd__xnor2_4 _19050_ (.A(_12332_),
    .B(_12336_),
    .Y(_12337_));
 sky130_fd_sc_hd__xnor2_1 _19051_ (.A(_12331_),
    .B(_12337_),
    .Y(_12338_));
 sky130_fd_sc_hd__nor2_1 _19052_ (.A(_12320_),
    .B(_12338_),
    .Y(_12339_));
 sky130_fd_sc_hd__and2_1 _19053_ (.A(_12320_),
    .B(_12338_),
    .X(_12340_));
 sky130_fd_sc_hd__nor2_1 _19054_ (.A(_12339_),
    .B(_12340_),
    .Y(_12341_));
 sky130_fd_sc_hd__nor3_1 _19055_ (.A(_12208_),
    .B(_12220_),
    .C(_12221_),
    .Y(_12342_));
 sky130_fd_sc_hd__buf_2 _19056_ (.A(_11712_),
    .X(_12343_));
 sky130_fd_sc_hd__nand2_1 _19057_ (.A(_11900_),
    .B(_12343_),
    .Y(_12344_));
 sky130_fd_sc_hd__and4_1 _19058_ (.A(_11904_),
    .B(_11110_),
    .C(_11054_),
    .D(_11170_),
    .X(_12345_));
 sky130_fd_sc_hd__a22o_1 _19059_ (.A1(_11905_),
    .A2(_11054_),
    .B1(_12098_),
    .B2(_11904_),
    .X(_12346_));
 sky130_fd_sc_hd__and2b_1 _19060_ (.A_N(_12345_),
    .B(_12346_),
    .X(_12347_));
 sky130_fd_sc_hd__xnor2_1 _19061_ (.A(_12344_),
    .B(_12347_),
    .Y(_12348_));
 sky130_fd_sc_hd__nand2_1 _19062_ (.A(_11268_),
    .B(_11134_),
    .Y(_12349_));
 sky130_fd_sc_hd__and4_1 _19063_ (.A(_11047_),
    .B(_10918_),
    .C(_11240_),
    .D(_11910_),
    .X(_12350_));
 sky130_fd_sc_hd__a22oi_2 _19064_ (.A1(_11903_),
    .A2(_11235_),
    .B1(_11455_),
    .B2(_11174_),
    .Y(_12351_));
 sky130_fd_sc_hd__or3_1 _19065_ (.A(_12349_),
    .B(_12350_),
    .C(_12351_),
    .X(_12352_));
 sky130_fd_sc_hd__o21ai_1 _19066_ (.A1(_12350_),
    .A2(_12351_),
    .B1(_12349_),
    .Y(_12353_));
 sky130_fd_sc_hd__o21bai_1 _19067_ (.A1(_12199_),
    .A2(_12201_),
    .B1_N(_12200_),
    .Y(_12354_));
 sky130_fd_sc_hd__and3_1 _19068_ (.A(_12352_),
    .B(_12353_),
    .C(_12354_),
    .X(_12355_));
 sky130_fd_sc_hd__a21o_1 _19069_ (.A1(_12352_),
    .A2(_12353_),
    .B1(_12354_),
    .X(_12356_));
 sky130_fd_sc_hd__and2b_1 _19070_ (.A_N(_12355_),
    .B(_12356_),
    .X(_12357_));
 sky130_fd_sc_hd__xnor2_1 _19071_ (.A(_12348_),
    .B(_12357_),
    .Y(_12358_));
 sky130_fd_sc_hd__or2b_1 _19072_ (.A(_12212_),
    .B_N(_12217_),
    .X(_12359_));
 sky130_fd_sc_hd__or2b_1 _19073_ (.A(_12211_),
    .B_N(_12218_),
    .X(_12360_));
 sky130_fd_sc_hd__clkbuf_4 _19074_ (.A(_10912_),
    .X(_12361_));
 sky130_fd_sc_hd__a31o_1 _19075_ (.A1(_12361_),
    .A2(_11444_),
    .A3(_12216_),
    .B1(_12214_),
    .X(_12362_));
 sky130_fd_sc_hd__o21bai_2 _19076_ (.A1(_12231_),
    .A2(_12236_),
    .B1_N(_12234_),
    .Y(_12363_));
 sky130_fd_sc_hd__clkbuf_2 _19077_ (.A(\genblk1.pcpi_mul.rs2[15] ),
    .X(_12364_));
 sky130_fd_sc_hd__nand2_1 _19078_ (.A(_10805_),
    .B(_12364_),
    .Y(_12365_));
 sky130_fd_sc_hd__nand4_2 _19079_ (.A(_10792_),
    .B(_10696_),
    .C(_11662_),
    .D(_11924_),
    .Y(_12366_));
 sky130_fd_sc_hd__a22o_1 _19080_ (.A1(_10848_),
    .A2(_11922_),
    .B1(_11924_),
    .B2(_10696_),
    .X(_12367_));
 sky130_fd_sc_hd__nand3b_1 _19081_ (.A_N(_12365_),
    .B(_12366_),
    .C(_12367_),
    .Y(_12368_));
 sky130_fd_sc_hd__a21bo_1 _19082_ (.A1(_12366_),
    .A2(_12367_),
    .B1_N(_12365_),
    .X(_12369_));
 sky130_fd_sc_hd__nand3_1 _19083_ (.A(_12363_),
    .B(_12368_),
    .C(_12369_),
    .Y(_12370_));
 sky130_fd_sc_hd__a21o_1 _19084_ (.A1(_12368_),
    .A2(_12369_),
    .B1(_12363_),
    .X(_12371_));
 sky130_fd_sc_hd__and3_1 _19085_ (.A(_12362_),
    .B(_12370_),
    .C(_12371_),
    .X(_12372_));
 sky130_fd_sc_hd__a21oi_1 _19086_ (.A1(_12370_),
    .A2(_12371_),
    .B1(_12362_),
    .Y(_12373_));
 sky130_fd_sc_hd__or2_1 _19087_ (.A(_12372_),
    .B(_12373_),
    .X(_12374_));
 sky130_fd_sc_hd__a21oi_2 _19088_ (.A1(_12359_),
    .A2(_12360_),
    .B1(_12374_),
    .Y(_12375_));
 sky130_fd_sc_hd__and3_1 _19089_ (.A(_12359_),
    .B(_12360_),
    .C(_12374_),
    .X(_12376_));
 sky130_fd_sc_hd__or3_2 _19090_ (.A(_12358_),
    .B(_12375_),
    .C(_12376_),
    .X(_12377_));
 sky130_fd_sc_hd__o21ai_1 _19091_ (.A1(_12375_),
    .A2(_12376_),
    .B1(_12358_),
    .Y(_12378_));
 sky130_fd_sc_hd__o211ai_2 _19092_ (.A1(_12220_),
    .A2(_12342_),
    .B1(_12377_),
    .C1(_12378_),
    .Y(_12379_));
 sky130_fd_sc_hd__a211o_1 _19093_ (.A1(_12377_),
    .A2(_12378_),
    .B1(_12220_),
    .C1(_12342_),
    .X(_12380_));
 sky130_fd_sc_hd__nand3_1 _19094_ (.A(_12341_),
    .B(_12379_),
    .C(_12380_),
    .Y(_12381_));
 sky130_fd_sc_hd__a21o_1 _19095_ (.A1(_12379_),
    .A2(_12380_),
    .B1(_12341_),
    .X(_12382_));
 sky130_fd_sc_hd__and3_1 _19096_ (.A(_12240_),
    .B(_12381_),
    .C(_12382_),
    .X(_12383_));
 sky130_fd_sc_hd__a21oi_1 _19097_ (.A1(_12381_),
    .A2(_12382_),
    .B1(_12240_),
    .Y(_12384_));
 sky130_fd_sc_hd__nor4_2 _19098_ (.A(_12318_),
    .B(_12319_),
    .C(_12383_),
    .D(_12384_),
    .Y(_12385_));
 sky130_fd_sc_hd__o22a_2 _19099_ (.A1(_12318_),
    .A2(_12319_),
    .B1(_12383_),
    .B2(_12384_),
    .X(_12386_));
 sky130_fd_sc_hd__a211oi_4 _19100_ (.A1(_12242_),
    .A2(_12244_),
    .B1(net342),
    .C1(_12386_),
    .Y(_12387_));
 sky130_fd_sc_hd__o211a_1 _19101_ (.A1(net342),
    .A2(_12386_),
    .B1(_12242_),
    .C1(_12244_),
    .X(_12388_));
 sky130_fd_sc_hd__or3_1 _19102_ (.A(_12265_),
    .B(_12387_),
    .C(_12388_),
    .X(_12389_));
 sky130_fd_sc_hd__o21ai_1 _19103_ (.A1(_12387_),
    .A2(_12388_),
    .B1(_12265_),
    .Y(_12390_));
 sky130_fd_sc_hd__o211a_1 _19104_ (.A1(_12246_),
    .A2(_12262_),
    .B1(_12389_),
    .C1(_12390_),
    .X(_12391_));
 sky130_fd_sc_hd__a211oi_1 _19105_ (.A1(_12389_),
    .A2(_12390_),
    .B1(_12246_),
    .C1(_12262_),
    .Y(_12392_));
 sky130_fd_sc_hd__nor3_1 _19106_ (.A(_12261_),
    .B(_12391_),
    .C(_12392_),
    .Y(_12393_));
 sky130_fd_sc_hd__o21a_1 _19107_ (.A1(_12391_),
    .A2(_12392_),
    .B1(_12261_),
    .X(_12394_));
 sky130_fd_sc_hd__or2_1 _19108_ (.A(_12393_),
    .B(_12394_),
    .X(_12395_));
 sky130_fd_sc_hd__or2b_1 _19109_ (.A(_12250_),
    .B_N(_12252_),
    .X(_12396_));
 sky130_fd_sc_hd__xnor2_1 _19110_ (.A(_12395_),
    .B(_12396_),
    .Y(_12397_));
 sky130_fd_sc_hd__and2b_1 _19111_ (.A_N(_12260_),
    .B(_12397_),
    .X(_12398_));
 sky130_fd_sc_hd__and2b_1 _19112_ (.A_N(_12397_),
    .B(_12260_),
    .X(_12399_));
 sky130_fd_sc_hd__nor2_1 _19113_ (.A(_12398_),
    .B(_12399_),
    .Y(_00068_));
 sky130_fd_sc_hd__or2_1 _19114_ (.A(_12263_),
    .B(_12264_),
    .X(_12400_));
 sky130_fd_sc_hd__nor3_1 _19115_ (.A(_12265_),
    .B(_12387_),
    .C(_12388_),
    .Y(_12401_));
 sky130_fd_sc_hd__nor2_1 _19116_ (.A(_12316_),
    .B(_12318_),
    .Y(_12402_));
 sky130_fd_sc_hd__nor2_1 _19117_ (.A(_12292_),
    .B(_12294_),
    .Y(_12403_));
 sky130_fd_sc_hd__xnor2_1 _19118_ (.A(_12402_),
    .B(_12403_),
    .Y(_12404_));
 sky130_fd_sc_hd__or2_1 _19119_ (.A(_12146_),
    .B(_12275_),
    .X(_12405_));
 sky130_fd_sc_hd__a211o_1 _19120_ (.A1(_12148_),
    .A2(_12272_),
    .B1(_12279_),
    .C1(_12276_),
    .X(_12406_));
 sky130_fd_sc_hd__or2b_1 _19121_ (.A(_12289_),
    .B_N(_12288_),
    .X(_12407_));
 sky130_fd_sc_hd__nand2_1 _19122_ (.A(_12280_),
    .B(_12290_),
    .Y(_12408_));
 sky130_fd_sc_hd__nand2_1 _19123_ (.A(_10640_),
    .B(_12282_),
    .Y(_12409_));
 sky130_fd_sc_hd__nand2_1 _19124_ (.A(_10740_),
    .B(_12282_),
    .Y(_12410_));
 sky130_fd_sc_hd__nor2_1 _19125_ (.A(_12272_),
    .B(_12410_),
    .Y(_12411_));
 sky130_fd_sc_hd__a21oi_1 _19126_ (.A1(_12275_),
    .A2(_12409_),
    .B1(_12411_),
    .Y(_12412_));
 sky130_fd_sc_hd__buf_2 _19127_ (.A(_12145_),
    .X(_12413_));
 sky130_fd_sc_hd__nand2_2 _19128_ (.A(_10625_),
    .B(_12413_),
    .Y(_12414_));
 sky130_fd_sc_hd__xnor2_1 _19129_ (.A(_12412_),
    .B(_12414_),
    .Y(_12415_));
 sky130_fd_sc_hd__clkbuf_4 _19130_ (.A(\genblk1.pcpi_mul.rs1[23] ),
    .X(_12416_));
 sky130_fd_sc_hd__nand2_1 _19131_ (.A(_10583_),
    .B(_12416_),
    .Y(_12417_));
 sky130_fd_sc_hd__and4_1 _19132_ (.A(_10661_),
    .B(_10707_),
    .C(_11829_),
    .D(_12069_),
    .X(_12418_));
 sky130_fd_sc_hd__a22oi_2 _19133_ (.A1(_11711_),
    .A2(_11946_),
    .B1(_11958_),
    .B2(_11710_),
    .Y(_12419_));
 sky130_fd_sc_hd__nor2_1 _19134_ (.A(_12418_),
    .B(_12419_),
    .Y(_12420_));
 sky130_fd_sc_hd__xnor2_1 _19135_ (.A(_12417_),
    .B(_12420_),
    .Y(_12421_));
 sky130_fd_sc_hd__o21ba_1 _19136_ (.A1(_12283_),
    .A2(_12286_),
    .B1_N(_12284_),
    .X(_12422_));
 sky130_fd_sc_hd__xnor2_1 _19137_ (.A(_12421_),
    .B(_12422_),
    .Y(_12423_));
 sky130_fd_sc_hd__xnor2_1 _19138_ (.A(_12415_),
    .B(_12423_),
    .Y(_12424_));
 sky130_fd_sc_hd__a21oi_1 _19139_ (.A1(_12407_),
    .A2(_12408_),
    .B1(_12424_),
    .Y(_12425_));
 sky130_fd_sc_hd__and3_1 _19140_ (.A(_12407_),
    .B(_12408_),
    .C(_12424_),
    .X(_12426_));
 sky130_fd_sc_hd__a211oi_1 _19141_ (.A1(_12405_),
    .A2(_12406_),
    .B1(_12425_),
    .C1(_12426_),
    .Y(_12427_));
 sky130_fd_sc_hd__o211a_1 _19142_ (.A1(_12425_),
    .A2(_12426_),
    .B1(_12405_),
    .C1(_12406_),
    .X(_12428_));
 sky130_fd_sc_hd__nand3_1 _19143_ (.A(_12296_),
    .B(_12306_),
    .C(_12307_),
    .Y(_12429_));
 sky130_fd_sc_hd__a21o_1 _19144_ (.A1(_12348_),
    .A2(_12356_),
    .B1(_12355_),
    .X(_12430_));
 sky130_fd_sc_hd__nand2_1 _19145_ (.A(_12300_),
    .B(_12302_),
    .Y(_12431_));
 sky130_fd_sc_hd__a31o_1 _19146_ (.A1(_10892_),
    .A2(_11277_),
    .A3(_12346_),
    .B1(_12345_),
    .X(_12432_));
 sky130_fd_sc_hd__nand4_2 _19147_ (.A(_10782_),
    .B(_11200_),
    .C(_11589_),
    .D(_12081_),
    .Y(_12433_));
 sky130_fd_sc_hd__a22o_1 _19148_ (.A1(_11085_),
    .A2(_11589_),
    .B1(_11597_),
    .B2(_12172_),
    .X(_12434_));
 sky130_fd_sc_hd__nand4_2 _19149_ (.A(_11508_),
    .B(_11708_),
    .C(_12433_),
    .D(_12434_),
    .Y(_12435_));
 sky130_fd_sc_hd__a22o_1 _19150_ (.A1(_10736_),
    .A2(_11819_),
    .B1(_12433_),
    .B2(_12434_),
    .X(_12436_));
 sky130_fd_sc_hd__nand3_2 _19151_ (.A(_12432_),
    .B(_12435_),
    .C(_12436_),
    .Y(_12437_));
 sky130_fd_sc_hd__a21o_1 _19152_ (.A1(_12435_),
    .A2(_12436_),
    .B1(_12432_),
    .X(_12438_));
 sky130_fd_sc_hd__nand3_2 _19153_ (.A(_12431_),
    .B(_12437_),
    .C(_12438_),
    .Y(_12439_));
 sky130_fd_sc_hd__a21o_1 _19154_ (.A1(_12437_),
    .A2(_12438_),
    .B1(_12431_),
    .X(_12440_));
 sky130_fd_sc_hd__and3_1 _19155_ (.A(_12430_),
    .B(_12439_),
    .C(_12440_),
    .X(_12441_));
 sky130_fd_sc_hd__a21oi_1 _19156_ (.A1(_12439_),
    .A2(_12440_),
    .B1(_12430_),
    .Y(_12442_));
 sky130_fd_sc_hd__a211oi_2 _19157_ (.A1(_12304_),
    .A2(_12306_),
    .B1(_12441_),
    .C1(_12442_),
    .Y(_12443_));
 sky130_fd_sc_hd__o211a_1 _19158_ (.A1(_12441_),
    .A2(_12442_),
    .B1(_12304_),
    .C1(_12306_),
    .X(_12444_));
 sky130_fd_sc_hd__a211oi_1 _19159_ (.A1(_12429_),
    .A2(_12310_),
    .B1(_12443_),
    .C1(_12444_),
    .Y(_12445_));
 sky130_fd_sc_hd__o211a_1 _19160_ (.A1(_12443_),
    .A2(_12444_),
    .B1(_12429_),
    .C1(_12310_),
    .X(_12446_));
 sky130_fd_sc_hd__or4_1 _19161_ (.A(_12427_),
    .B(_12428_),
    .C(_12445_),
    .D(_12446_),
    .X(_12447_));
 sky130_fd_sc_hd__o22ai_1 _19162_ (.A1(_12427_),
    .A2(_12428_),
    .B1(_12445_),
    .B2(_12446_),
    .Y(_12448_));
 sky130_fd_sc_hd__and3b_1 _19163_ (.A_N(_12379_),
    .B(_12447_),
    .C(_12448_),
    .X(_12449_));
 sky130_fd_sc_hd__a21boi_1 _19164_ (.A1(_12447_),
    .A2(_12448_),
    .B1_N(_12379_),
    .Y(_12450_));
 sky130_fd_sc_hd__a211oi_1 _19165_ (.A1(_12312_),
    .A2(_12314_),
    .B1(_12449_),
    .C1(_12450_),
    .Y(_12451_));
 sky130_fd_sc_hd__o211a_1 _19166_ (.A1(_12449_),
    .A2(_12450_),
    .B1(_12312_),
    .C1(_12314_),
    .X(_12452_));
 sky130_fd_sc_hd__nand2_1 _19167_ (.A(_12331_),
    .B(_12337_),
    .Y(_12453_));
 sky130_fd_sc_hd__nand2_1 _19168_ (.A(_10855_),
    .B(_11770_),
    .Y(_12454_));
 sky130_fd_sc_hd__and4_1 _19169_ (.A(_10800_),
    .B(_10718_),
    .C(_12333_),
    .D(_12232_),
    .X(_12455_));
 sky130_fd_sc_hd__a22o_1 _19170_ (.A1(_10664_),
    .A2(_12333_),
    .B1(_12020_),
    .B2(_10800_),
    .X(_12456_));
 sky130_fd_sc_hd__and2b_1 _19171_ (.A_N(_12455_),
    .B(_12456_),
    .X(_12457_));
 sky130_fd_sc_hd__xnor2_2 _19172_ (.A(_12454_),
    .B(_12457_),
    .Y(_12458_));
 sky130_vsdinv _19173_ (.A(_12458_),
    .Y(_12459_));
 sky130_fd_sc_hd__buf_2 _19174_ (.A(\genblk1.pcpi_mul.rs2[21] ),
    .X(_12460_));
 sky130_fd_sc_hd__nand2_2 _19175_ (.A(_11777_),
    .B(_12460_),
    .Y(_12461_));
 sky130_fd_sc_hd__buf_1 _19176_ (.A(\genblk1.pcpi_mul.rs2[23] ),
    .X(_12462_));
 sky130_fd_sc_hd__and4_1 _19177_ (.A(_10709_),
    .B(_10704_),
    .C(_12321_),
    .D(_12462_),
    .X(_12463_));
 sky130_fd_sc_hd__clkbuf_2 _19178_ (.A(\genblk1.pcpi_mul.rs2[23] ),
    .X(_12464_));
 sky130_fd_sc_hd__a22o_1 _19179_ (.A1(_10704_),
    .A2(_12321_),
    .B1(_12464_),
    .B2(_10709_),
    .X(_12465_));
 sky130_fd_sc_hd__and2b_1 _19180_ (.A_N(_12463_),
    .B(_12465_),
    .X(_12466_));
 sky130_fd_sc_hd__xnor2_4 _19181_ (.A(_12461_),
    .B(_12466_),
    .Y(_12467_));
 sky130_fd_sc_hd__xnor2_1 _19182_ (.A(_12330_),
    .B(_12467_),
    .Y(_12468_));
 sky130_fd_sc_hd__xnor2_1 _19183_ (.A(_12459_),
    .B(_12468_),
    .Y(_12469_));
 sky130_fd_sc_hd__nor2_1 _19184_ (.A(_12453_),
    .B(_12469_),
    .Y(_12470_));
 sky130_fd_sc_hd__and2_1 _19185_ (.A(_12453_),
    .B(_12469_),
    .X(_12471_));
 sky130_fd_sc_hd__or2_1 _19186_ (.A(_12470_),
    .B(_12471_),
    .X(_12472_));
 sky130_vsdinv _19187_ (.A(_12375_),
    .Y(_12473_));
 sky130_fd_sc_hd__nand2_1 _19188_ (.A(_11190_),
    .B(_11482_),
    .Y(_12474_));
 sky130_fd_sc_hd__and4_1 _19189_ (.A(_11141_),
    .B(_11144_),
    .C(_11260_),
    .D(_11371_),
    .X(_12475_));
 sky130_fd_sc_hd__a22o_1 _19190_ (.A1(_11144_),
    .A2(_11260_),
    .B1(_11276_),
    .B2(_11141_),
    .X(_12476_));
 sky130_fd_sc_hd__and2b_1 _19191_ (.A_N(_12475_),
    .B(_12476_),
    .X(_12477_));
 sky130_fd_sc_hd__xnor2_2 _19192_ (.A(_12474_),
    .B(_12477_),
    .Y(_12478_));
 sky130_fd_sc_hd__nand2_1 _19193_ (.A(_11159_),
    .B(_11134_),
    .Y(_12479_));
 sky130_fd_sc_hd__and4_1 _19194_ (.A(_10918_),
    .B(_11154_),
    .C(_11234_),
    .D(_11457_),
    .X(_12480_));
 sky130_fd_sc_hd__a22oi_2 _19195_ (.A1(_10976_),
    .A2(_11795_),
    .B1(_11455_),
    .B2(_11903_),
    .Y(_12481_));
 sky130_fd_sc_hd__or3_1 _19196_ (.A(_12479_),
    .B(_12480_),
    .C(_12481_),
    .X(_12482_));
 sky130_fd_sc_hd__o21ai_1 _19197_ (.A1(_12480_),
    .A2(_12481_),
    .B1(_12479_),
    .Y(_12483_));
 sky130_fd_sc_hd__o21bai_1 _19198_ (.A1(_12349_),
    .A2(_12351_),
    .B1_N(_12350_),
    .Y(_12484_));
 sky130_fd_sc_hd__and3_1 _19199_ (.A(_12482_),
    .B(_12483_),
    .C(_12484_),
    .X(_12485_));
 sky130_fd_sc_hd__a21o_1 _19200_ (.A1(_12482_),
    .A2(_12483_),
    .B1(_12484_),
    .X(_12486_));
 sky130_fd_sc_hd__and2b_1 _19201_ (.A_N(_12485_),
    .B(_12486_),
    .X(_12487_));
 sky130_fd_sc_hd__xnor2_1 _19202_ (.A(_12478_),
    .B(_12487_),
    .Y(_12488_));
 sky130_fd_sc_hd__nand2_2 _19203_ (.A(_12366_),
    .B(_12368_),
    .Y(_12489_));
 sky130_fd_sc_hd__a31o_1 _19204_ (.A1(_10665_),
    .A2(_11769_),
    .A3(_12335_),
    .B1(_12334_),
    .X(_12490_));
 sky130_fd_sc_hd__nand4_2 _19205_ (.A(_10978_),
    .B(_10849_),
    .C(_11554_),
    .D(_11780_),
    .Y(_12491_));
 sky130_fd_sc_hd__a22o_1 _19206_ (.A1(_10851_),
    .A2(_11661_),
    .B1(_11657_),
    .B2(_10756_),
    .X(_12492_));
 sky130_fd_sc_hd__nand4_2 _19207_ (.A(_11048_),
    .B(_11443_),
    .C(_12491_),
    .D(_12492_),
    .Y(_12493_));
 sky130_fd_sc_hd__a22o_1 _19208_ (.A1(_10967_),
    .A2(_11443_),
    .B1(_12491_),
    .B2(_12492_),
    .X(_12494_));
 sky130_fd_sc_hd__nand3_2 _19209_ (.A(_12490_),
    .B(_12493_),
    .C(_12494_),
    .Y(_12495_));
 sky130_fd_sc_hd__a21o_1 _19210_ (.A1(_12493_),
    .A2(_12494_),
    .B1(_12490_),
    .X(_12496_));
 sky130_fd_sc_hd__nand3_1 _19211_ (.A(_12489_),
    .B(_12495_),
    .C(_12496_),
    .Y(_12497_));
 sky130_fd_sc_hd__a21o_1 _19212_ (.A1(_12495_),
    .A2(_12496_),
    .B1(_12489_),
    .X(_12498_));
 sky130_fd_sc_hd__a21bo_1 _19213_ (.A1(_12362_),
    .A2(_12371_),
    .B1_N(_12370_),
    .X(_12499_));
 sky130_fd_sc_hd__and3_1 _19214_ (.A(_12497_),
    .B(_12498_),
    .C(_12499_),
    .X(_12500_));
 sky130_fd_sc_hd__a21oi_1 _19215_ (.A1(_12497_),
    .A2(_12498_),
    .B1(_12499_),
    .Y(_12501_));
 sky130_fd_sc_hd__or3_2 _19216_ (.A(_12488_),
    .B(_12500_),
    .C(_12501_),
    .X(_12502_));
 sky130_fd_sc_hd__o21ai_1 _19217_ (.A1(_12500_),
    .A2(_12501_),
    .B1(_12488_),
    .Y(_12503_));
 sky130_fd_sc_hd__and3_1 _19218_ (.A(_12339_),
    .B(_12502_),
    .C(_12503_),
    .X(_12504_));
 sky130_fd_sc_hd__a21oi_1 _19219_ (.A1(_12502_),
    .A2(_12503_),
    .B1(_12339_),
    .Y(_12505_));
 sky130_fd_sc_hd__a211oi_2 _19220_ (.A1(_12473_),
    .A2(_12377_),
    .B1(_12504_),
    .C1(_12505_),
    .Y(_12506_));
 sky130_fd_sc_hd__o211a_1 _19221_ (.A1(_12504_),
    .A2(_12505_),
    .B1(_12473_),
    .C1(_12377_),
    .X(_12507_));
 sky130_fd_sc_hd__or3_2 _19222_ (.A(_12472_),
    .B(_12506_),
    .C(_12507_),
    .X(_12508_));
 sky130_fd_sc_hd__o21ai_1 _19223_ (.A1(_12506_),
    .A2(_12507_),
    .B1(_12472_),
    .Y(_12509_));
 sky130_fd_sc_hd__nand3b_2 _19224_ (.A_N(_12381_),
    .B(_12508_),
    .C(_12509_),
    .Y(_12510_));
 sky130_fd_sc_hd__a21bo_1 _19225_ (.A1(_12508_),
    .A2(_12509_),
    .B1_N(_12381_),
    .X(_12511_));
 sky130_fd_sc_hd__or4bb_2 _19226_ (.A(_12451_),
    .B(_12452_),
    .C_N(_12510_),
    .D_N(_12511_),
    .X(_12512_));
 sky130_fd_sc_hd__a2bb2o_1 _19227_ (.A1_N(_12451_),
    .A2_N(_12452_),
    .B1(_12510_),
    .B2(_12511_),
    .X(_12513_));
 sky130_fd_sc_hd__o211a_1 _19228_ (.A1(_12383_),
    .A2(_12385_),
    .B1(_12512_),
    .C1(_12513_),
    .X(_12514_));
 sky130_fd_sc_hd__a211oi_2 _19229_ (.A1(_12512_),
    .A2(_12513_),
    .B1(_12383_),
    .C1(_12385_),
    .Y(_12515_));
 sky130_fd_sc_hd__or3_2 _19230_ (.A(_12404_),
    .B(_12514_),
    .C(_12515_),
    .X(_12516_));
 sky130_fd_sc_hd__o21ai_2 _19231_ (.A1(_12514_),
    .A2(_12515_),
    .B1(_12404_),
    .Y(_12517_));
 sky130_fd_sc_hd__o211a_1 _19232_ (.A1(_12387_),
    .A2(_12401_),
    .B1(_12516_),
    .C1(_12517_),
    .X(_12518_));
 sky130_fd_sc_hd__a211oi_2 _19233_ (.A1(_12516_),
    .A2(_12517_),
    .B1(_12387_),
    .C1(_12401_),
    .Y(_12519_));
 sky130_fd_sc_hd__or3_2 _19234_ (.A(_12400_),
    .B(_12518_),
    .C(_12519_),
    .X(_12520_));
 sky130_fd_sc_hd__o21ai_2 _19235_ (.A1(_12518_),
    .A2(_12519_),
    .B1(_12400_),
    .Y(_12521_));
 sky130_fd_sc_hd__a211oi_2 _19236_ (.A1(_12520_),
    .A2(_12521_),
    .B1(_12391_),
    .C1(_12393_),
    .Y(_12522_));
 sky130_fd_sc_hd__o211a_1 _19237_ (.A1(_12391_),
    .A2(_12393_),
    .B1(_12520_),
    .C1(_12521_),
    .X(_12523_));
 sky130_fd_sc_hd__nor2_1 _19238_ (.A(_12522_),
    .B(_12523_),
    .Y(_12524_));
 sky130_fd_sc_hd__and2b_1 _19239_ (.A_N(_12395_),
    .B(_12396_),
    .X(_12525_));
 sky130_fd_sc_hd__nor2_1 _19240_ (.A(_12525_),
    .B(_12398_),
    .Y(_12526_));
 sky130_fd_sc_hd__xnor2_1 _19241_ (.A(_12524_),
    .B(_12526_),
    .Y(_00069_));
 sky130_fd_sc_hd__or2_1 _19242_ (.A(_12402_),
    .B(_12403_),
    .X(_12527_));
 sky130_fd_sc_hd__nor3_1 _19243_ (.A(_12404_),
    .B(_12514_),
    .C(_12515_),
    .Y(_12528_));
 sky130_fd_sc_hd__nor2_1 _19244_ (.A(_12449_),
    .B(_12451_),
    .Y(_12529_));
 sky130_fd_sc_hd__nor2_1 _19245_ (.A(_12425_),
    .B(_12427_),
    .Y(_12530_));
 sky130_fd_sc_hd__xnor2_1 _19246_ (.A(_12529_),
    .B(_12530_),
    .Y(_12531_));
 sky130_fd_sc_hd__or2b_1 _19247_ (.A(_12445_),
    .B_N(_12447_),
    .X(_12532_));
 sky130_fd_sc_hd__or2_1 _19248_ (.A(_12272_),
    .B(_12410_),
    .X(_12533_));
 sky130_fd_sc_hd__a211o_1 _19249_ (.A1(_12275_),
    .A2(_12409_),
    .B1(_12414_),
    .C1(_12411_),
    .X(_12534_));
 sky130_fd_sc_hd__or2b_1 _19250_ (.A(_12422_),
    .B_N(_12421_),
    .X(_12535_));
 sky130_fd_sc_hd__nand2_1 _19251_ (.A(_12415_),
    .B(_12423_),
    .Y(_12536_));
 sky130_fd_sc_hd__clkbuf_4 _19252_ (.A(\genblk1.pcpi_mul.rs1[23] ),
    .X(_12537_));
 sky130_fd_sc_hd__buf_4 _19253_ (.A(_12537_),
    .X(_12538_));
 sky130_fd_sc_hd__nand2_2 _19254_ (.A(_10747_),
    .B(_12538_),
    .Y(_12539_));
 sky130_fd_sc_hd__nand2_2 _19255_ (.A(_10611_),
    .B(_12416_),
    .Y(_12540_));
 sky130_fd_sc_hd__nor2_1 _19256_ (.A(_12409_),
    .B(_12540_),
    .Y(_12541_));
 sky130_fd_sc_hd__a21oi_1 _19257_ (.A1(_12410_),
    .A2(_12539_),
    .B1(_12541_),
    .Y(_12542_));
 sky130_fd_sc_hd__clkbuf_4 _19258_ (.A(_12154_),
    .X(_12543_));
 sky130_fd_sc_hd__nand2_2 _19259_ (.A(_11704_),
    .B(_12543_),
    .Y(_12544_));
 sky130_fd_sc_hd__xnor2_1 _19260_ (.A(_12542_),
    .B(_12544_),
    .Y(_12545_));
 sky130_fd_sc_hd__clkbuf_4 _19261_ (.A(\genblk1.pcpi_mul.rs1[24] ),
    .X(_12546_));
 sky130_fd_sc_hd__nand2_1 _19262_ (.A(_10583_),
    .B(_12546_),
    .Y(_12547_));
 sky130_fd_sc_hd__and4_1 _19263_ (.A(_10700_),
    .B(_10803_),
    .C(_12069_),
    .D(_12078_),
    .X(_12548_));
 sky130_fd_sc_hd__a22oi_2 _19264_ (.A1(_11711_),
    .A2(_11958_),
    .B1(_12147_),
    .B2(_10671_),
    .Y(_12549_));
 sky130_fd_sc_hd__nor2_1 _19265_ (.A(_12548_),
    .B(_12549_),
    .Y(_12550_));
 sky130_fd_sc_hd__xnor2_1 _19266_ (.A(_12547_),
    .B(_12550_),
    .Y(_12551_));
 sky130_fd_sc_hd__o21ba_1 _19267_ (.A1(_12417_),
    .A2(_12419_),
    .B1_N(_12418_),
    .X(_12552_));
 sky130_fd_sc_hd__xnor2_1 _19268_ (.A(_12551_),
    .B(_12552_),
    .Y(_12553_));
 sky130_fd_sc_hd__xnor2_1 _19269_ (.A(_12545_),
    .B(_12553_),
    .Y(_12554_));
 sky130_fd_sc_hd__a21oi_1 _19270_ (.A1(_12535_),
    .A2(_12536_),
    .B1(_12554_),
    .Y(_12555_));
 sky130_fd_sc_hd__and3_1 _19271_ (.A(_12535_),
    .B(_12536_),
    .C(_12554_),
    .X(_12556_));
 sky130_fd_sc_hd__a211oi_1 _19272_ (.A1(_12533_),
    .A2(_12534_),
    .B1(_12555_),
    .C1(_12556_),
    .Y(_12557_));
 sky130_fd_sc_hd__o211a_1 _19273_ (.A1(_12555_),
    .A2(_12556_),
    .B1(_12533_),
    .C1(_12534_),
    .X(_12558_));
 sky130_fd_sc_hd__a21o_1 _19274_ (.A1(_12478_),
    .A2(_12486_),
    .B1(_12485_),
    .X(_12559_));
 sky130_fd_sc_hd__nand2_1 _19275_ (.A(_12433_),
    .B(_12435_),
    .Y(_12560_));
 sky130_fd_sc_hd__clkbuf_4 _19276_ (.A(_11476_),
    .X(_12561_));
 sky130_fd_sc_hd__a31o_1 _19277_ (.A1(_11900_),
    .A2(_12561_),
    .A3(_12476_),
    .B1(_12475_),
    .X(_12562_));
 sky130_fd_sc_hd__nand2_1 _19278_ (.A(_10787_),
    .B(_11830_),
    .Y(_12563_));
 sky130_fd_sc_hd__nand4_2 _19279_ (.A(_11082_),
    .B(_10998_),
    .C(_11698_),
    .D(_11707_),
    .Y(_12564_));
 sky130_fd_sc_hd__a22o_1 _19280_ (.A1(_10998_),
    .A2(_12081_),
    .B1(_11707_),
    .B2(_10782_),
    .X(_12565_));
 sky130_fd_sc_hd__nand3b_1 _19281_ (.A_N(_12563_),
    .B(_12564_),
    .C(_12565_),
    .Y(_12566_));
 sky130_fd_sc_hd__a21bo_1 _19282_ (.A1(_12564_),
    .A2(_12565_),
    .B1_N(_12563_),
    .X(_12567_));
 sky130_fd_sc_hd__nand3_2 _19283_ (.A(_12562_),
    .B(_12566_),
    .C(_12567_),
    .Y(_12568_));
 sky130_fd_sc_hd__a21o_1 _19284_ (.A1(_12566_),
    .A2(_12567_),
    .B1(_12562_),
    .X(_12569_));
 sky130_fd_sc_hd__nand3_2 _19285_ (.A(_12560_),
    .B(_12568_),
    .C(_12569_),
    .Y(_12570_));
 sky130_fd_sc_hd__a21o_1 _19286_ (.A1(_12568_),
    .A2(_12569_),
    .B1(_12560_),
    .X(_12571_));
 sky130_fd_sc_hd__and3_1 _19287_ (.A(_12559_),
    .B(_12570_),
    .C(_12571_),
    .X(_12572_));
 sky130_fd_sc_hd__a21oi_1 _19288_ (.A1(_12570_),
    .A2(_12571_),
    .B1(_12559_),
    .Y(_12573_));
 sky130_fd_sc_hd__a211o_1 _19289_ (.A1(_12437_),
    .A2(_12439_),
    .B1(_12572_),
    .C1(_12573_),
    .X(_12574_));
 sky130_fd_sc_hd__o211ai_1 _19290_ (.A1(_12572_),
    .A2(_12573_),
    .B1(_12437_),
    .C1(_12439_),
    .Y(_12575_));
 sky130_fd_sc_hd__o211ai_1 _19291_ (.A1(_12441_),
    .A2(_12443_),
    .B1(_12574_),
    .C1(_12575_),
    .Y(_12576_));
 sky130_fd_sc_hd__a211o_1 _19292_ (.A1(_12574_),
    .A2(_12575_),
    .B1(_12441_),
    .C1(_12443_),
    .X(_12577_));
 sky130_fd_sc_hd__or4bb_1 _19293_ (.A(_12557_),
    .B(_12558_),
    .C_N(_12576_),
    .D_N(_12577_),
    .X(_12578_));
 sky130_fd_sc_hd__a2bb2o_1 _19294_ (.A1_N(_12557_),
    .A2_N(_12558_),
    .B1(_12576_),
    .B2(_12577_),
    .X(_12579_));
 sky130_fd_sc_hd__o211ai_1 _19295_ (.A1(_12504_),
    .A2(_12506_),
    .B1(_12578_),
    .C1(_12579_),
    .Y(_12580_));
 sky130_fd_sc_hd__a211o_1 _19296_ (.A1(_12578_),
    .A2(_12579_),
    .B1(_12504_),
    .C1(_12506_),
    .X(_12581_));
 sky130_fd_sc_hd__and3_1 _19297_ (.A(_12532_),
    .B(_12580_),
    .C(_12581_),
    .X(_12582_));
 sky130_fd_sc_hd__a21oi_1 _19298_ (.A1(_12580_),
    .A2(_12581_),
    .B1(_12532_),
    .Y(_12583_));
 sky130_fd_sc_hd__buf_2 _19299_ (.A(\genblk1.pcpi_mul.rs2[24] ),
    .X(_12584_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19300_ (.A(_12584_),
    .X(_12585_));
 sky130_fd_sc_hd__clkbuf_4 _19301_ (.A(_12585_),
    .X(_12586_));
 sky130_fd_sc_hd__clkbuf_4 _19302_ (.A(_12586_),
    .X(_12587_));
 sky130_fd_sc_hd__nand2_2 _19303_ (.A(_10591_),
    .B(_12587_),
    .Y(_12588_));
 sky130_fd_sc_hd__nand2_1 _19304_ (.A(_12330_),
    .B(_12467_),
    .Y(_12589_));
 sky130_fd_sc_hd__or2_1 _19305_ (.A(_12459_),
    .B(_12468_),
    .X(_12590_));
 sky130_fd_sc_hd__clkbuf_4 _19306_ (.A(_11894_),
    .X(_12591_));
 sky130_fd_sc_hd__nand2_2 _19307_ (.A(_11404_),
    .B(_12591_),
    .Y(_12592_));
 sky130_fd_sc_hd__buf_1 _19308_ (.A(\genblk1.pcpi_mul.rs2[19] ),
    .X(_12593_));
 sky130_fd_sc_hd__and4_1 _19309_ (.A(_10718_),
    .B(\genblk1.pcpi_mul.rs1[5] ),
    .C(_12593_),
    .D(\genblk1.pcpi_mul.rs2[20] ),
    .X(_12594_));
 sky130_fd_sc_hd__a22o_1 _19310_ (.A1(_10793_),
    .A2(_12593_),
    .B1(_12232_),
    .B2(_10718_),
    .X(_12595_));
 sky130_fd_sc_hd__and2b_1 _19311_ (.A_N(_12594_),
    .B(_12595_),
    .X(_12596_));
 sky130_fd_sc_hd__xnor2_2 _19312_ (.A(_12592_),
    .B(_12596_),
    .Y(_12597_));
 sky130_fd_sc_hd__nand2_1 _19313_ (.A(_10675_),
    .B(_12460_),
    .Y(_12598_));
 sky130_fd_sc_hd__and4_1 _19314_ (.A(_10634_),
    .B(_10752_),
    .C(_12327_),
    .D(_12464_),
    .X(_12599_));
 sky130_fd_sc_hd__buf_2 _19315_ (.A(_12462_),
    .X(_12600_));
 sky130_fd_sc_hd__a22oi_2 _19316_ (.A1(_10754_),
    .A2(_12322_),
    .B1(_12600_),
    .B2(_10594_),
    .Y(_12601_));
 sky130_fd_sc_hd__nor2_1 _19317_ (.A(_12599_),
    .B(_12601_),
    .Y(_12602_));
 sky130_fd_sc_hd__xnor2_2 _19318_ (.A(_12598_),
    .B(_12602_),
    .Y(_12603_));
 sky130_fd_sc_hd__a31o_1 _19319_ (.A1(_10608_),
    .A2(_12226_),
    .A3(_12465_),
    .B1(_12463_),
    .X(_12604_));
 sky130_fd_sc_hd__xor2_1 _19320_ (.A(_12603_),
    .B(_12604_),
    .X(_12605_));
 sky130_fd_sc_hd__xnor2_1 _19321_ (.A(_12597_),
    .B(_12605_),
    .Y(_12606_));
 sky130_fd_sc_hd__a21oi_2 _19322_ (.A1(_12589_),
    .A2(_12590_),
    .B1(_12606_),
    .Y(_12607_));
 sky130_fd_sc_hd__and3_1 _19323_ (.A(_12589_),
    .B(_12590_),
    .C(_12606_),
    .X(_12608_));
 sky130_fd_sc_hd__or3_1 _19324_ (.A(_12588_),
    .B(_12607_),
    .C(_12608_),
    .X(_12609_));
 sky130_fd_sc_hd__o21ai_1 _19325_ (.A1(_12607_),
    .A2(_12608_),
    .B1(_12588_),
    .Y(_12610_));
 sky130_fd_sc_hd__and2_1 _19326_ (.A(_12609_),
    .B(_12610_),
    .X(_12611_));
 sky130_fd_sc_hd__nand3_1 _19327_ (.A(_12497_),
    .B(_12498_),
    .C(_12499_),
    .Y(_12612_));
 sky130_fd_sc_hd__nand2_1 _19328_ (.A(_10960_),
    .B(_11961_),
    .Y(_12613_));
 sky130_fd_sc_hd__and4_1 _19329_ (.A(_10955_),
    .B(_11143_),
    .C(_11275_),
    .D(_11379_),
    .X(_12614_));
 sky130_fd_sc_hd__a22o_1 _19330_ (.A1(_11106_),
    .A2(_11275_),
    .B1(_11379_),
    .B2(_10955_),
    .X(_12615_));
 sky130_fd_sc_hd__and2b_1 _19331_ (.A_N(_12614_),
    .B(_12615_),
    .X(_12616_));
 sky130_fd_sc_hd__xnor2_1 _19332_ (.A(_12613_),
    .B(_12616_),
    .Y(_12617_));
 sky130_fd_sc_hd__nand2_1 _19333_ (.A(_11349_),
    .B(_11170_),
    .Y(_12618_));
 sky130_fd_sc_hd__and4_1 _19334_ (.A(\genblk1.pcpi_mul.rs1[10] ),
    .B(\genblk1.pcpi_mul.rs1[11] ),
    .C(_11239_),
    .D(_11457_),
    .X(_12619_));
 sky130_fd_sc_hd__a22oi_2 _19335_ (.A1(_11066_),
    .A2(_11234_),
    .B1(_11910_),
    .B2(_11154_),
    .Y(_12620_));
 sky130_fd_sc_hd__or3_1 _19336_ (.A(_12618_),
    .B(_12619_),
    .C(_12620_),
    .X(_12621_));
 sky130_fd_sc_hd__o21ai_1 _19337_ (.A1(_12619_),
    .A2(_12620_),
    .B1(_12618_),
    .Y(_12622_));
 sky130_fd_sc_hd__o21bai_1 _19338_ (.A1(_12479_),
    .A2(_12481_),
    .B1_N(_12480_),
    .Y(_12623_));
 sky130_fd_sc_hd__and3_1 _19339_ (.A(_12621_),
    .B(_12622_),
    .C(_12623_),
    .X(_12624_));
 sky130_fd_sc_hd__a21o_1 _19340_ (.A1(_12621_),
    .A2(_12622_),
    .B1(_12623_),
    .X(_12625_));
 sky130_fd_sc_hd__and2b_1 _19341_ (.A_N(_12624_),
    .B(_12625_),
    .X(_12626_));
 sky130_fd_sc_hd__xnor2_1 _19342_ (.A(_12617_),
    .B(_12626_),
    .Y(_12627_));
 sky130_fd_sc_hd__nand2_2 _19343_ (.A(_12491_),
    .B(_12493_),
    .Y(_12628_));
 sky130_fd_sc_hd__a31o_1 _19344_ (.A1(_10790_),
    .A2(_11769_),
    .A3(_12456_),
    .B1(_12455_),
    .X(_12629_));
 sky130_fd_sc_hd__nand2_1 _19345_ (.A(_11903_),
    .B(_12364_),
    .Y(_12630_));
 sky130_fd_sc_hd__nand4_2 _19346_ (.A(_10849_),
    .B(_11047_),
    .C(_11554_),
    .D(_11780_),
    .Y(_12631_));
 sky130_fd_sc_hd__a22o_1 _19347_ (.A1(_10907_),
    .A2(_11554_),
    .B1(_11657_),
    .B2(_10851_),
    .X(_12632_));
 sky130_fd_sc_hd__nand3b_1 _19348_ (.A_N(_12630_),
    .B(_12631_),
    .C(_12632_),
    .Y(_12633_));
 sky130_fd_sc_hd__a21bo_1 _19349_ (.A1(_12631_),
    .A2(_12632_),
    .B1_N(_12630_),
    .X(_12634_));
 sky130_fd_sc_hd__nand3_1 _19350_ (.A(_12629_),
    .B(_12633_),
    .C(_12634_),
    .Y(_12635_));
 sky130_fd_sc_hd__a21o_1 _19351_ (.A1(_12633_),
    .A2(_12634_),
    .B1(_12629_),
    .X(_12636_));
 sky130_fd_sc_hd__nand3_1 _19352_ (.A(_12628_),
    .B(_12635_),
    .C(_12636_),
    .Y(_12637_));
 sky130_fd_sc_hd__a21o_1 _19353_ (.A1(_12635_),
    .A2(_12636_),
    .B1(_12628_),
    .X(_12638_));
 sky130_fd_sc_hd__a21bo_1 _19354_ (.A1(_12489_),
    .A2(_12496_),
    .B1_N(_12495_),
    .X(_12639_));
 sky130_fd_sc_hd__and3_1 _19355_ (.A(_12637_),
    .B(_12638_),
    .C(_12639_),
    .X(_12640_));
 sky130_fd_sc_hd__a21oi_1 _19356_ (.A1(_12637_),
    .A2(_12638_),
    .B1(_12639_),
    .Y(_12641_));
 sky130_fd_sc_hd__or3_1 _19357_ (.A(_12627_),
    .B(_12640_),
    .C(_12641_),
    .X(_12642_));
 sky130_fd_sc_hd__clkbuf_2 _19358_ (.A(_12642_),
    .X(_12643_));
 sky130_fd_sc_hd__o21ai_1 _19359_ (.A1(_12640_),
    .A2(_12641_),
    .B1(_12627_),
    .Y(_12644_));
 sky130_fd_sc_hd__and3_1 _19360_ (.A(_12470_),
    .B(_12643_),
    .C(_12644_),
    .X(_12645_));
 sky130_fd_sc_hd__a21oi_1 _19361_ (.A1(_12643_),
    .A2(_12644_),
    .B1(_12470_),
    .Y(_12646_));
 sky130_fd_sc_hd__a211o_1 _19362_ (.A1(_12612_),
    .A2(_12502_),
    .B1(_12645_),
    .C1(_12646_),
    .X(_12647_));
 sky130_fd_sc_hd__o211ai_1 _19363_ (.A1(_12645_),
    .A2(_12646_),
    .B1(_12612_),
    .C1(_12502_),
    .Y(_12648_));
 sky130_fd_sc_hd__and3_1 _19364_ (.A(_12611_),
    .B(_12647_),
    .C(_12648_),
    .X(_12649_));
 sky130_fd_sc_hd__a21oi_1 _19365_ (.A1(_12647_),
    .A2(_12648_),
    .B1(_12611_),
    .Y(_12650_));
 sky130_fd_sc_hd__nor3_1 _19366_ (.A(_12508_),
    .B(_12649_),
    .C(_12650_),
    .Y(_12651_));
 sky130_fd_sc_hd__o21a_1 _19367_ (.A1(_12649_),
    .A2(_12650_),
    .B1(_12508_),
    .X(_12652_));
 sky130_fd_sc_hd__nor4_1 _19368_ (.A(_12582_),
    .B(_12583_),
    .C(net347),
    .D(_12652_),
    .Y(_12653_));
 sky130_fd_sc_hd__o22a_1 _19369_ (.A1(_12582_),
    .A2(_12583_),
    .B1(net347),
    .B2(_12652_),
    .X(_12654_));
 sky130_fd_sc_hd__a211oi_2 _19370_ (.A1(_12510_),
    .A2(_12512_),
    .B1(net341),
    .C1(_12654_),
    .Y(_12655_));
 sky130_fd_sc_hd__o211a_1 _19371_ (.A1(net341),
    .A2(_12654_),
    .B1(_12510_),
    .C1(_12512_),
    .X(_12656_));
 sky130_fd_sc_hd__or3_1 _19372_ (.A(_12531_),
    .B(_12655_),
    .C(_12656_),
    .X(_12657_));
 sky130_fd_sc_hd__o21ai_1 _19373_ (.A1(_12655_),
    .A2(_12656_),
    .B1(_12531_),
    .Y(_12658_));
 sky130_fd_sc_hd__o211a_1 _19374_ (.A1(_12514_),
    .A2(_12528_),
    .B1(_12657_),
    .C1(_12658_),
    .X(_12659_));
 sky130_fd_sc_hd__a211oi_1 _19375_ (.A1(_12657_),
    .A2(_12658_),
    .B1(_12514_),
    .C1(_12528_),
    .Y(_12660_));
 sky130_fd_sc_hd__or3_1 _19376_ (.A(_12527_),
    .B(_12659_),
    .C(_12660_),
    .X(_12661_));
 sky130_fd_sc_hd__o21ai_1 _19377_ (.A1(_12659_),
    .A2(_12660_),
    .B1(_12527_),
    .Y(_12662_));
 sky130_fd_sc_hd__o21bai_2 _19378_ (.A1(_12400_),
    .A2(_12519_),
    .B1_N(_12518_),
    .Y(_12663_));
 sky130_fd_sc_hd__and3_1 _19379_ (.A(_12661_),
    .B(_12662_),
    .C(_12663_),
    .X(_12664_));
 sky130_fd_sc_hd__a21oi_1 _19380_ (.A1(_12661_),
    .A2(_12662_),
    .B1(_12663_),
    .Y(_12665_));
 sky130_fd_sc_hd__or2_1 _19381_ (.A(_12664_),
    .B(_12665_),
    .X(_12666_));
 sky130_fd_sc_hd__nand4b_1 _19382_ (.A_N(_12130_),
    .B(_12256_),
    .C(_12397_),
    .D(_12524_),
    .Y(_12667_));
 sky130_fd_sc_hd__a211o_1 _19383_ (.A1(_11542_),
    .A2(_11547_),
    .B1(_12131_),
    .C1(_12667_),
    .X(_12668_));
 sky130_fd_sc_hd__and4b_1 _19384_ (.A_N(_12130_),
    .B(_12256_),
    .C(_12397_),
    .D(_12524_),
    .X(_12669_));
 sky130_fd_sc_hd__and3_1 _19385_ (.A(_12397_),
    .B(_12259_),
    .C(_12524_),
    .X(_12670_));
 sky130_vsdinv _19386_ (.A(_12522_),
    .Y(_12671_));
 sky130_fd_sc_hd__a21o_1 _19387_ (.A1(_12525_),
    .A2(_12671_),
    .B1(_12523_),
    .X(_12672_));
 sky130_fd_sc_hd__a211oi_2 _19388_ (.A1(_12133_),
    .A2(_12669_),
    .B1(_12670_),
    .C1(_12672_),
    .Y(_12673_));
 sky130_fd_sc_hd__and2_2 _19389_ (.A(_12668_),
    .B(_12673_),
    .X(_12674_));
 sky130_fd_sc_hd__xor2_1 _19390_ (.A(_12666_),
    .B(_12674_),
    .X(_00070_));
 sky130_fd_sc_hd__or2_1 _19391_ (.A(_12529_),
    .B(_12530_),
    .X(_12675_));
 sky130_fd_sc_hd__nor3_1 _19392_ (.A(_12531_),
    .B(_12655_),
    .C(_12656_),
    .Y(_12676_));
 sky130_fd_sc_hd__a21boi_1 _19393_ (.A1(_12532_),
    .A2(_12581_),
    .B1_N(_12580_),
    .Y(_12677_));
 sky130_fd_sc_hd__nor2_1 _19394_ (.A(_12555_),
    .B(_12557_),
    .Y(_12678_));
 sky130_fd_sc_hd__or2_1 _19395_ (.A(_12677_),
    .B(_12678_),
    .X(_12679_));
 sky130_fd_sc_hd__nand2_1 _19396_ (.A(_12677_),
    .B(_12678_),
    .Y(_12680_));
 sky130_fd_sc_hd__nand2_1 _19397_ (.A(_12679_),
    .B(_12680_),
    .Y(_12681_));
 sky130_fd_sc_hd__nand2_1 _19398_ (.A(_12576_),
    .B(_12578_),
    .Y(_12682_));
 sky130_fd_sc_hd__nand3_1 _19399_ (.A(_12470_),
    .B(_12643_),
    .C(_12644_),
    .Y(_12683_));
 sky130_fd_sc_hd__or2_1 _19400_ (.A(_12409_),
    .B(_12540_),
    .X(_12684_));
 sky130_fd_sc_hd__a211o_1 _19401_ (.A1(_12410_),
    .A2(_12539_),
    .B1(_12544_),
    .C1(_12541_),
    .X(_12685_));
 sky130_fd_sc_hd__or2b_1 _19402_ (.A(_12552_),
    .B_N(_12551_),
    .X(_12686_));
 sky130_fd_sc_hd__nand2_1 _19403_ (.A(_12545_),
    .B(_12553_),
    .Y(_12687_));
 sky130_fd_sc_hd__clkbuf_4 _19404_ (.A(\genblk1.pcpi_mul.rs1[24] ),
    .X(_12688_));
 sky130_fd_sc_hd__nand2_1 _19405_ (.A(_10639_),
    .B(_12688_),
    .Y(_12689_));
 sky130_fd_sc_hd__buf_4 _19406_ (.A(\genblk1.pcpi_mul.rs1[24] ),
    .X(_12690_));
 sky130_fd_sc_hd__nand2_1 _19407_ (.A(_10740_),
    .B(_12690_),
    .Y(_12691_));
 sky130_fd_sc_hd__nor2_1 _19408_ (.A(_12539_),
    .B(_12691_),
    .Y(_12692_));
 sky130_fd_sc_hd__a21oi_1 _19409_ (.A1(_12540_),
    .A2(_12689_),
    .B1(_12692_),
    .Y(_12693_));
 sky130_fd_sc_hd__buf_2 _19410_ (.A(_12282_),
    .X(_12694_));
 sky130_fd_sc_hd__nand2_2 _19411_ (.A(_10625_),
    .B(_12694_),
    .Y(_12695_));
 sky130_fd_sc_hd__xnor2_1 _19412_ (.A(_12693_),
    .B(_12695_),
    .Y(_12696_));
 sky130_fd_sc_hd__and4_1 _19413_ (.A(_10670_),
    .B(_10916_),
    .C(_12143_),
    .D(_12153_),
    .X(_12697_));
 sky130_fd_sc_hd__a22oi_4 _19414_ (.A1(_10803_),
    .A2(_12078_),
    .B1(_12273_),
    .B2(_10700_),
    .Y(_12698_));
 sky130_fd_sc_hd__nor2_1 _19415_ (.A(_12697_),
    .B(_12698_),
    .Y(_12699_));
 sky130_fd_sc_hd__buf_2 _19416_ (.A(\genblk1.pcpi_mul.rs1[25] ),
    .X(_12700_));
 sky130_fd_sc_hd__nand2_1 _19417_ (.A(_10695_),
    .B(_12700_),
    .Y(_12701_));
 sky130_fd_sc_hd__xnor2_1 _19418_ (.A(_12699_),
    .B(_12701_),
    .Y(_12702_));
 sky130_fd_sc_hd__o21ba_1 _19419_ (.A1(_12547_),
    .A2(_12549_),
    .B1_N(_12548_),
    .X(_12703_));
 sky130_fd_sc_hd__xnor2_1 _19420_ (.A(_12702_),
    .B(_12703_),
    .Y(_12704_));
 sky130_fd_sc_hd__xnor2_1 _19421_ (.A(_12696_),
    .B(_12704_),
    .Y(_12705_));
 sky130_fd_sc_hd__a21oi_1 _19422_ (.A1(_12686_),
    .A2(_12687_),
    .B1(_12705_),
    .Y(_12706_));
 sky130_fd_sc_hd__and3_1 _19423_ (.A(_12686_),
    .B(_12687_),
    .C(_12705_),
    .X(_12707_));
 sky130_fd_sc_hd__a211oi_1 _19424_ (.A1(_12684_),
    .A2(_12685_),
    .B1(_12706_),
    .C1(_12707_),
    .Y(_12708_));
 sky130_fd_sc_hd__o211a_1 _19425_ (.A1(_12706_),
    .A2(_12707_),
    .B1(_12684_),
    .C1(_12685_),
    .X(_12709_));
 sky130_fd_sc_hd__nand3_1 _19426_ (.A(_12559_),
    .B(_12570_),
    .C(_12571_),
    .Y(_12710_));
 sky130_fd_sc_hd__a21o_1 _19427_ (.A1(_12617_),
    .A2(_12625_),
    .B1(_12624_),
    .X(_12711_));
 sky130_fd_sc_hd__nand2_1 _19428_ (.A(_12564_),
    .B(_12566_),
    .Y(_12712_));
 sky130_fd_sc_hd__a31o_1 _19429_ (.A1(_11189_),
    .A2(_11489_),
    .A3(_12615_),
    .B1(_12614_),
    .X(_12713_));
 sky130_fd_sc_hd__clkbuf_2 _19430_ (.A(\genblk1.pcpi_mul.rs1[17] ),
    .X(_12714_));
 sky130_fd_sc_hd__nand4_2 _19431_ (.A(_12172_),
    .B(_11195_),
    .C(_12714_),
    .D(_11829_),
    .Y(_12715_));
 sky130_fd_sc_hd__a22o_1 _19432_ (.A1(_10837_),
    .A2(_12714_),
    .B1(_11945_),
    .B2(_10995_),
    .X(_12716_));
 sky130_fd_sc_hd__nand4_2 _19433_ (.A(_10993_),
    .B(_12067_),
    .C(_12715_),
    .D(_12716_),
    .Y(_12717_));
 sky130_fd_sc_hd__a22o_1 _19434_ (.A1(_10787_),
    .A2(_11958_),
    .B1(_12715_),
    .B2(_12716_),
    .X(_12718_));
 sky130_fd_sc_hd__nand3_2 _19435_ (.A(_12713_),
    .B(_12717_),
    .C(_12718_),
    .Y(_12719_));
 sky130_fd_sc_hd__a21o_1 _19436_ (.A1(_12717_),
    .A2(_12718_),
    .B1(_12713_),
    .X(_12720_));
 sky130_fd_sc_hd__nand3_2 _19437_ (.A(_12712_),
    .B(_12719_),
    .C(_12720_),
    .Y(_12721_));
 sky130_fd_sc_hd__a21o_1 _19438_ (.A1(_12719_),
    .A2(_12720_),
    .B1(_12712_),
    .X(_12722_));
 sky130_fd_sc_hd__and3_2 _19439_ (.A(_12711_),
    .B(_12721_),
    .C(_12722_),
    .X(_12723_));
 sky130_fd_sc_hd__a21oi_2 _19440_ (.A1(_12721_),
    .A2(_12722_),
    .B1(_12711_),
    .Y(_12724_));
 sky130_fd_sc_hd__a211oi_4 _19441_ (.A1(_12568_),
    .A2(_12570_),
    .B1(_12723_),
    .C1(_12724_),
    .Y(_12725_));
 sky130_fd_sc_hd__o211a_1 _19442_ (.A1(_12723_),
    .A2(_12724_),
    .B1(_12568_),
    .C1(_12570_),
    .X(_12726_));
 sky130_fd_sc_hd__a211oi_2 _19443_ (.A1(_12710_),
    .A2(_12574_),
    .B1(_12725_),
    .C1(_12726_),
    .Y(_12727_));
 sky130_fd_sc_hd__o211a_1 _19444_ (.A1(_12725_),
    .A2(_12726_),
    .B1(_12710_),
    .C1(_12574_),
    .X(_12728_));
 sky130_fd_sc_hd__nor4_1 _19445_ (.A(_12708_),
    .B(_12709_),
    .C(_12727_),
    .D(_12728_),
    .Y(_12729_));
 sky130_fd_sc_hd__o22a_1 _19446_ (.A1(_12708_),
    .A2(_12709_),
    .B1(_12727_),
    .B2(_12728_),
    .X(_12730_));
 sky130_fd_sc_hd__a211o_1 _19447_ (.A1(_12683_),
    .A2(_12647_),
    .B1(net365),
    .C1(_12730_),
    .X(_12731_));
 sky130_fd_sc_hd__o211ai_2 _19448_ (.A1(net365),
    .A2(_12730_),
    .B1(_12683_),
    .C1(_12647_),
    .Y(_12732_));
 sky130_fd_sc_hd__nand3_2 _19449_ (.A(_12682_),
    .B(_12731_),
    .C(_12732_),
    .Y(_12733_));
 sky130_fd_sc_hd__a21o_1 _19450_ (.A1(_12731_),
    .A2(_12732_),
    .B1(_12682_),
    .X(_12734_));
 sky130_fd_sc_hd__nand3_1 _19451_ (.A(_12637_),
    .B(_12638_),
    .C(_12639_),
    .Y(_12735_));
 sky130_fd_sc_hd__nand2_1 _19452_ (.A(_11189_),
    .B(_11598_),
    .Y(_12736_));
 sky130_fd_sc_hd__and4_1 _19453_ (.A(_11140_),
    .B(_11143_),
    .C(_11480_),
    .D(_11588_),
    .X(_12737_));
 sky130_fd_sc_hd__a22o_1 _19454_ (.A1(_11143_),
    .A2(_11480_),
    .B1(_11588_),
    .B2(_11140_),
    .X(_12738_));
 sky130_fd_sc_hd__and2b_1 _19455_ (.A_N(_12737_),
    .B(_12738_),
    .X(_12739_));
 sky130_fd_sc_hd__xnor2_1 _19456_ (.A(_12736_),
    .B(_12739_),
    .Y(_12740_));
 sky130_fd_sc_hd__nand2_1 _19457_ (.A(_11349_),
    .B(_11275_),
    .Y(_12741_));
 sky130_fd_sc_hd__and4_1 _19458_ (.A(\genblk1.pcpi_mul.rs1[11] ),
    .B(\genblk1.pcpi_mul.rs1[12] ),
    .C(_11239_),
    .D(_11352_),
    .X(_12742_));
 sky130_fd_sc_hd__a22oi_2 _19459_ (.A1(_11170_),
    .A2(_11234_),
    .B1(_11910_),
    .B2(_11066_),
    .Y(_12743_));
 sky130_fd_sc_hd__or3_1 _19460_ (.A(_12741_),
    .B(_12742_),
    .C(_12743_),
    .X(_12744_));
 sky130_fd_sc_hd__o21ai_1 _19461_ (.A1(_12742_),
    .A2(_12743_),
    .B1(_12741_),
    .Y(_12745_));
 sky130_fd_sc_hd__o21bai_1 _19462_ (.A1(_12618_),
    .A2(_12620_),
    .B1_N(_12619_),
    .Y(_12746_));
 sky130_fd_sc_hd__and3_1 _19463_ (.A(_12744_),
    .B(_12745_),
    .C(_12746_),
    .X(_12747_));
 sky130_fd_sc_hd__a21o_1 _19464_ (.A1(_12744_),
    .A2(_12745_),
    .B1(_12746_),
    .X(_12748_));
 sky130_fd_sc_hd__and2b_1 _19465_ (.A_N(_12747_),
    .B(_12748_),
    .X(_12749_));
 sky130_fd_sc_hd__xnor2_1 _19466_ (.A(_12740_),
    .B(_12749_),
    .Y(_12750_));
 sky130_fd_sc_hd__nand2_1 _19467_ (.A(_12631_),
    .B(_12633_),
    .Y(_12751_));
 sky130_fd_sc_hd__a31o_1 _19468_ (.A1(_10792_),
    .A2(_11769_),
    .A3(_12595_),
    .B1(_12594_),
    .X(_12752_));
 sky130_fd_sc_hd__nand4_2 _19469_ (.A(_10907_),
    .B(_10918_),
    .C(_11554_),
    .D(_11657_),
    .Y(_12753_));
 sky130_fd_sc_hd__a22o_1 _19470_ (.A1(_10918_),
    .A2(_11661_),
    .B1(\genblk1.pcpi_mul.rs2[17] ),
    .B2(\genblk1.pcpi_mul.rs1[8] ),
    .X(_12754_));
 sky130_fd_sc_hd__nand4_2 _19471_ (.A(_11155_),
    .B(_11443_),
    .C(_12753_),
    .D(_12754_),
    .Y(_12755_));
 sky130_fd_sc_hd__a22o_1 _19472_ (.A1(_11268_),
    .A2(_12364_),
    .B1(_12753_),
    .B2(_12754_),
    .X(_12756_));
 sky130_fd_sc_hd__nand3_1 _19473_ (.A(_12752_),
    .B(_12755_),
    .C(_12756_),
    .Y(_12757_));
 sky130_fd_sc_hd__a21o_1 _19474_ (.A1(_12755_),
    .A2(_12756_),
    .B1(_12752_),
    .X(_12758_));
 sky130_fd_sc_hd__nand3_1 _19475_ (.A(_12751_),
    .B(_12757_),
    .C(_12758_),
    .Y(_12759_));
 sky130_fd_sc_hd__a21o_1 _19476_ (.A1(_12757_),
    .A2(_12758_),
    .B1(_12751_),
    .X(_12760_));
 sky130_fd_sc_hd__a21bo_1 _19477_ (.A1(_12628_),
    .A2(_12636_),
    .B1_N(_12635_),
    .X(_12761_));
 sky130_fd_sc_hd__and3_1 _19478_ (.A(_12759_),
    .B(_12760_),
    .C(_12761_),
    .X(_12762_));
 sky130_fd_sc_hd__a21oi_1 _19479_ (.A1(_12759_),
    .A2(_12760_),
    .B1(_12761_),
    .Y(_12763_));
 sky130_fd_sc_hd__or3_2 _19480_ (.A(_12750_),
    .B(_12762_),
    .C(_12763_),
    .X(_12764_));
 sky130_fd_sc_hd__o21ai_1 _19481_ (.A1(_12762_),
    .A2(_12763_),
    .B1(_12750_),
    .Y(_12765_));
 sky130_fd_sc_hd__and3_2 _19482_ (.A(_12607_),
    .B(_12764_),
    .C(_12765_),
    .X(_12766_));
 sky130_fd_sc_hd__a21oi_1 _19483_ (.A1(_12764_),
    .A2(_12765_),
    .B1(_12607_),
    .Y(_12767_));
 sky130_fd_sc_hd__a211o_1 _19484_ (.A1(_12735_),
    .A2(_12643_),
    .B1(_12766_),
    .C1(_12767_),
    .X(_12768_));
 sky130_fd_sc_hd__o211ai_2 _19485_ (.A1(_12766_),
    .A2(_12767_),
    .B1(_12735_),
    .C1(_12643_),
    .Y(_12769_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19486_ (.A(\genblk1.pcpi_mul.rs2[25] ),
    .X(_12770_));
 sky130_fd_sc_hd__buf_2 _19487_ (.A(_12770_),
    .X(_12771_));
 sky130_fd_sc_hd__clkbuf_4 _19488_ (.A(_12771_),
    .X(_12772_));
 sky130_fd_sc_hd__buf_4 _19489_ (.A(_12772_),
    .X(_12773_));
 sky130_fd_sc_hd__a22oi_4 _19490_ (.A1(_10597_),
    .A2(_12587_),
    .B1(_12773_),
    .B2(_10590_),
    .Y(_12774_));
 sky130_fd_sc_hd__clkbuf_2 _19491_ (.A(\genblk1.pcpi_mul.rs2[24] ),
    .X(_12775_));
 sky130_fd_sc_hd__buf_2 _19492_ (.A(_12770_),
    .X(_12776_));
 sky130_fd_sc_hd__and4_1 _19493_ (.A(_10588_),
    .B(_10635_),
    .C(_12775_),
    .D(_12776_),
    .X(_12777_));
 sky130_fd_sc_hd__nor2_2 _19494_ (.A(_12774_),
    .B(_12777_),
    .Y(_12778_));
 sky130_fd_sc_hd__and2_1 _19495_ (.A(_12603_),
    .B(_12604_),
    .X(_12779_));
 sky130_fd_sc_hd__a21oi_2 _19496_ (.A1(_12597_),
    .A2(_12605_),
    .B1(_12779_),
    .Y(_12780_));
 sky130_fd_sc_hd__nand2_1 _19497_ (.A(_11405_),
    .B(_11895_),
    .Y(_12781_));
 sky130_fd_sc_hd__and4_1 _19498_ (.A(\genblk1.pcpi_mul.rs1[6] ),
    .B(\genblk1.pcpi_mul.rs1[5] ),
    .C(_12593_),
    .D(\genblk1.pcpi_mul.rs2[20] ),
    .X(_12782_));
 sky130_fd_sc_hd__a22o_1 _19499_ (.A1(_10756_),
    .A2(_12593_),
    .B1(\genblk1.pcpi_mul.rs2[20] ),
    .B2(\genblk1.pcpi_mul.rs1[5] ),
    .X(_12783_));
 sky130_fd_sc_hd__and2b_1 _19500_ (.A_N(_12782_),
    .B(_12783_),
    .X(_12784_));
 sky130_fd_sc_hd__xnor2_2 _19501_ (.A(_12781_),
    .B(_12784_),
    .Y(_12785_));
 sky130_fd_sc_hd__nand2_2 _19502_ (.A(_10744_),
    .B(_12460_),
    .Y(_12786_));
 sky130_fd_sc_hd__and4_1 _19503_ (.A(\genblk1.pcpi_mul.rs1[2] ),
    .B(_10647_),
    .C(_12321_),
    .D(_12462_),
    .X(_12787_));
 sky130_fd_sc_hd__a22o_1 _19504_ (.A1(_10647_),
    .A2(_12321_),
    .B1(_12462_),
    .B2(_10606_),
    .X(_12788_));
 sky130_fd_sc_hd__and2b_1 _19505_ (.A_N(_12787_),
    .B(_12788_),
    .X(_12789_));
 sky130_fd_sc_hd__xnor2_4 _19506_ (.A(_12786_),
    .B(_12789_),
    .Y(_12790_));
 sky130_fd_sc_hd__o21ba_2 _19507_ (.A1(_12598_),
    .A2(_12601_),
    .B1_N(_12599_),
    .X(_12791_));
 sky130_fd_sc_hd__xnor2_2 _19508_ (.A(_12790_),
    .B(_12791_),
    .Y(_12792_));
 sky130_fd_sc_hd__xnor2_2 _19509_ (.A(_12785_),
    .B(_12792_),
    .Y(_12793_));
 sky130_fd_sc_hd__xor2_2 _19510_ (.A(_12780_),
    .B(_12793_),
    .X(_12794_));
 sky130_fd_sc_hd__xnor2_2 _19511_ (.A(_12778_),
    .B(_12794_),
    .Y(_12795_));
 sky130_fd_sc_hd__xor2_1 _19512_ (.A(_12609_),
    .B(_12795_),
    .X(_12796_));
 sky130_fd_sc_hd__nand3_2 _19513_ (.A(_12768_),
    .B(_12769_),
    .C(_12796_),
    .Y(_12797_));
 sky130_fd_sc_hd__a21o_1 _19514_ (.A1(_12768_),
    .A2(_12769_),
    .B1(_12796_),
    .X(_12798_));
 sky130_fd_sc_hd__nand3_2 _19515_ (.A(_12649_),
    .B(_12797_),
    .C(_12798_),
    .Y(_12799_));
 sky130_fd_sc_hd__a21o_1 _19516_ (.A1(_12797_),
    .A2(_12798_),
    .B1(_12649_),
    .X(_12800_));
 sky130_fd_sc_hd__nand4_2 _19517_ (.A(_12733_),
    .B(_12734_),
    .C(_12799_),
    .D(_12800_),
    .Y(_12801_));
 sky130_fd_sc_hd__a22o_1 _19518_ (.A1(_12733_),
    .A2(_12734_),
    .B1(_12799_),
    .B2(_12800_),
    .X(_12802_));
 sky130_fd_sc_hd__o211a_1 _19519_ (.A1(_12651_),
    .A2(net416),
    .B1(_12801_),
    .C1(_12802_),
    .X(_12803_));
 sky130_fd_sc_hd__a211oi_1 _19520_ (.A1(_12801_),
    .A2(_12802_),
    .B1(_12651_),
    .C1(net416),
    .Y(_12804_));
 sky130_fd_sc_hd__or3_1 _19521_ (.A(_12681_),
    .B(_12803_),
    .C(_12804_),
    .X(_12805_));
 sky130_fd_sc_hd__o21ai_1 _19522_ (.A1(_12803_),
    .A2(_12804_),
    .B1(_12681_),
    .Y(_12806_));
 sky130_fd_sc_hd__o211a_1 _19523_ (.A1(_12655_),
    .A2(_12676_),
    .B1(_12805_),
    .C1(_12806_),
    .X(_12807_));
 sky130_fd_sc_hd__a211oi_1 _19524_ (.A1(_12805_),
    .A2(_12806_),
    .B1(_12655_),
    .C1(_12676_),
    .Y(_12808_));
 sky130_fd_sc_hd__or3_1 _19525_ (.A(_12675_),
    .B(_12807_),
    .C(_12808_),
    .X(_12809_));
 sky130_fd_sc_hd__o21ai_1 _19526_ (.A1(_12807_),
    .A2(_12808_),
    .B1(_12675_),
    .Y(_12810_));
 sky130_fd_sc_hd__nor3_1 _19527_ (.A(_12527_),
    .B(_12659_),
    .C(_12660_),
    .Y(_12811_));
 sky130_fd_sc_hd__a211oi_2 _19528_ (.A1(_12809_),
    .A2(_12810_),
    .B1(_12659_),
    .C1(_12811_),
    .Y(_12812_));
 sky130_fd_sc_hd__o211ai_1 _19529_ (.A1(_12659_),
    .A2(_12811_),
    .B1(_12809_),
    .C1(_12810_),
    .Y(_12813_));
 sky130_fd_sc_hd__and2b_1 _19530_ (.A_N(_12812_),
    .B(_12813_),
    .X(_12814_));
 sky130_fd_sc_hd__o21ba_1 _19531_ (.A1(_12666_),
    .A2(_12674_),
    .B1_N(_12664_),
    .X(_12815_));
 sky130_fd_sc_hd__xnor2_1 _19532_ (.A(_12814_),
    .B(_12815_),
    .Y(_00071_));
 sky130_fd_sc_hd__nor3_1 _19533_ (.A(_12675_),
    .B(_12807_),
    .C(_12808_),
    .Y(_12816_));
 sky130_fd_sc_hd__nor3_1 _19534_ (.A(_12681_),
    .B(_12803_),
    .C(_12804_),
    .Y(_12817_));
 sky130_fd_sc_hd__nand2_1 _19535_ (.A(_12731_),
    .B(_12733_),
    .Y(_12818_));
 sky130_fd_sc_hd__nor2_1 _19536_ (.A(_12706_),
    .B(_12708_),
    .Y(_12819_));
 sky130_fd_sc_hd__xor2_1 _19537_ (.A(_12818_),
    .B(_12819_),
    .X(_12820_));
 sky130_fd_sc_hd__a211oi_1 _19538_ (.A1(_12735_),
    .A2(_12643_),
    .B1(_12766_),
    .C1(_12767_),
    .Y(_12821_));
 sky130_fd_sc_hd__or2_1 _19539_ (.A(_12539_),
    .B(_12691_),
    .X(_12822_));
 sky130_fd_sc_hd__a211o_1 _19540_ (.A1(_12540_),
    .A2(_12689_),
    .B1(_12695_),
    .C1(_12692_),
    .X(_12823_));
 sky130_fd_sc_hd__or2b_1 _19541_ (.A(_12703_),
    .B_N(_12702_),
    .X(_12824_));
 sky130_fd_sc_hd__nand2_1 _19542_ (.A(_12696_),
    .B(_12704_),
    .Y(_12825_));
 sky130_fd_sc_hd__nand2_1 _19543_ (.A(_10747_),
    .B(_12700_),
    .Y(_12826_));
 sky130_fd_sc_hd__nand2_1 _19544_ (.A(_10610_),
    .B(_12700_),
    .Y(_12827_));
 sky130_fd_sc_hd__nor2_1 _19545_ (.A(_12689_),
    .B(_12827_),
    .Y(_12828_));
 sky130_fd_sc_hd__a21oi_1 _19546_ (.A1(_12691_),
    .A2(_12826_),
    .B1(_12828_),
    .Y(_12829_));
 sky130_fd_sc_hd__clkbuf_4 _19547_ (.A(_12537_),
    .X(_12830_));
 sky130_fd_sc_hd__nand2_2 _19548_ (.A(_10624_),
    .B(_12830_),
    .Y(_12831_));
 sky130_fd_sc_hd__xnor2_1 _19549_ (.A(_12829_),
    .B(_12831_),
    .Y(_12832_));
 sky130_fd_sc_hd__nand2_1 _19550_ (.A(_10582_),
    .B(\genblk1.pcpi_mul.rs1[26] ),
    .Y(_12833_));
 sky130_fd_sc_hd__and4_1 _19551_ (.A(_10699_),
    .B(_10706_),
    .C(\genblk1.pcpi_mul.rs1[21] ),
    .D(\genblk1.pcpi_mul.rs1[22] ),
    .X(_12834_));
 sky130_fd_sc_hd__a22oi_2 _19552_ (.A1(_10916_),
    .A2(_12153_),
    .B1(_12281_),
    .B2(_10802_),
    .Y(_12835_));
 sky130_fd_sc_hd__nor2_1 _19553_ (.A(_12834_),
    .B(_12835_),
    .Y(_12836_));
 sky130_fd_sc_hd__xnor2_1 _19554_ (.A(_12833_),
    .B(_12836_),
    .Y(_12837_));
 sky130_fd_sc_hd__o21ba_1 _19555_ (.A1(_12698_),
    .A2(_12701_),
    .B1_N(_12697_),
    .X(_12838_));
 sky130_fd_sc_hd__xnor2_1 _19556_ (.A(_12837_),
    .B(_12838_),
    .Y(_12839_));
 sky130_fd_sc_hd__xnor2_1 _19557_ (.A(_12832_),
    .B(_12839_),
    .Y(_12840_));
 sky130_fd_sc_hd__a21oi_1 _19558_ (.A1(_12824_),
    .A2(_12825_),
    .B1(_12840_),
    .Y(_12841_));
 sky130_fd_sc_hd__and3_1 _19559_ (.A(_12824_),
    .B(_12825_),
    .C(_12840_),
    .X(_12842_));
 sky130_fd_sc_hd__a211oi_1 _19560_ (.A1(_12822_),
    .A2(_12823_),
    .B1(_12841_),
    .C1(_12842_),
    .Y(_12843_));
 sky130_fd_sc_hd__o211a_1 _19561_ (.A1(_12841_),
    .A2(_12842_),
    .B1(_12822_),
    .C1(_12823_),
    .X(_12844_));
 sky130_fd_sc_hd__a21o_1 _19562_ (.A1(_12740_),
    .A2(_12748_),
    .B1(_12747_),
    .X(_12845_));
 sky130_fd_sc_hd__nand2_1 _19563_ (.A(_12715_),
    .B(_12717_),
    .Y(_12846_));
 sky130_fd_sc_hd__a31o_1 _19564_ (.A1(_11189_),
    .A2(_12081_),
    .A3(_12738_),
    .B1(_12737_),
    .X(_12847_));
 sky130_fd_sc_hd__nand2_1 _19565_ (.A(_10735_),
    .B(_12143_),
    .Y(_12848_));
 sky130_fd_sc_hd__nand4_2 _19566_ (.A(_10995_),
    .B(_10837_),
    .C(_11945_),
    .D(_11957_),
    .Y(_12849_));
 sky130_fd_sc_hd__a22o_1 _19567_ (.A1(_10839_),
    .A2(_11945_),
    .B1(\genblk1.pcpi_mul.rs1[19] ),
    .B2(_10836_),
    .X(_12850_));
 sky130_fd_sc_hd__nand3b_2 _19568_ (.A_N(_12848_),
    .B(_12849_),
    .C(_12850_),
    .Y(_12851_));
 sky130_fd_sc_hd__a21bo_1 _19569_ (.A1(_12849_),
    .A2(_12850_),
    .B1_N(_12848_),
    .X(_12852_));
 sky130_fd_sc_hd__nand3_4 _19570_ (.A(_12847_),
    .B(_12851_),
    .C(_12852_),
    .Y(_12853_));
 sky130_fd_sc_hd__a21o_1 _19571_ (.A1(_12851_),
    .A2(_12852_),
    .B1(_12847_),
    .X(_12854_));
 sky130_fd_sc_hd__nand3_4 _19572_ (.A(_12846_),
    .B(_12853_),
    .C(_12854_),
    .Y(_12855_));
 sky130_fd_sc_hd__a21o_1 _19573_ (.A1(_12853_),
    .A2(_12854_),
    .B1(_12846_),
    .X(_12856_));
 sky130_fd_sc_hd__and3_1 _19574_ (.A(_12845_),
    .B(_12855_),
    .C(_12856_),
    .X(_12857_));
 sky130_fd_sc_hd__a21oi_1 _19575_ (.A1(_12855_),
    .A2(_12856_),
    .B1(_12845_),
    .Y(_12858_));
 sky130_fd_sc_hd__a211o_2 _19576_ (.A1(_12719_),
    .A2(_12721_),
    .B1(_12857_),
    .C1(_12858_),
    .X(_12859_));
 sky130_fd_sc_hd__o211ai_2 _19577_ (.A1(_12857_),
    .A2(_12858_),
    .B1(_12719_),
    .C1(_12721_),
    .Y(_12860_));
 sky130_fd_sc_hd__o211ai_4 _19578_ (.A1(_12723_),
    .A2(_12725_),
    .B1(_12859_),
    .C1(_12860_),
    .Y(_12861_));
 sky130_fd_sc_hd__a211o_1 _19579_ (.A1(_12859_),
    .A2(_12860_),
    .B1(_12723_),
    .C1(_12725_),
    .X(_12862_));
 sky130_fd_sc_hd__or4bb_2 _19580_ (.A(_12843_),
    .B(_12844_),
    .C_N(_12861_),
    .D_N(_12862_),
    .X(_12863_));
 sky130_fd_sc_hd__a2bb2o_1 _19581_ (.A1_N(_12843_),
    .A2_N(_12844_),
    .B1(_12861_),
    .B2(_12862_),
    .X(_12864_));
 sky130_fd_sc_hd__o211ai_2 _19582_ (.A1(_12766_),
    .A2(_12821_),
    .B1(_12863_),
    .C1(_12864_),
    .Y(_12865_));
 sky130_fd_sc_hd__a211o_1 _19583_ (.A1(_12863_),
    .A2(_12864_),
    .B1(_12766_),
    .C1(_12821_),
    .X(_12866_));
 sky130_fd_sc_hd__o211a_1 _19584_ (.A1(_12727_),
    .A2(net420),
    .B1(_12865_),
    .C1(_12866_),
    .X(_12867_));
 sky130_fd_sc_hd__a211oi_1 _19585_ (.A1(_12865_),
    .A2(_12866_),
    .B1(_12727_),
    .C1(net420),
    .Y(_12868_));
 sky130_fd_sc_hd__or2_1 _19586_ (.A(_12609_),
    .B(_12795_),
    .X(_12869_));
 sky130_fd_sc_hd__nand3_1 _19587_ (.A(_12759_),
    .B(_12760_),
    .C(_12761_),
    .Y(_12870_));
 sky130_fd_sc_hd__nor2_1 _19588_ (.A(_12780_),
    .B(_12793_),
    .Y(_12871_));
 sky130_fd_sc_hd__nand2_1 _19589_ (.A(_10892_),
    .B(_12074_),
    .Y(_12872_));
 sky130_fd_sc_hd__and4_1 _19590_ (.A(_10955_),
    .B(_11106_),
    .C(_11488_),
    .D(_11697_),
    .X(_12873_));
 sky130_fd_sc_hd__a22o_1 _19591_ (.A1(_11110_),
    .A2(_11488_),
    .B1(_11597_),
    .B2(_10962_),
    .X(_12874_));
 sky130_fd_sc_hd__and2b_1 _19592_ (.A_N(_12873_),
    .B(_12874_),
    .X(_12875_));
 sky130_fd_sc_hd__xnor2_1 _19593_ (.A(_12872_),
    .B(_12875_),
    .Y(_12876_));
 sky130_fd_sc_hd__nand2_1 _19594_ (.A(_11349_),
    .B(_11480_),
    .Y(_12877_));
 sky130_fd_sc_hd__and4_1 _19595_ (.A(\genblk1.pcpi_mul.rs1[12] ),
    .B(_11239_),
    .C(\genblk1.pcpi_mul.rs1[13] ),
    .D(_11352_),
    .X(_12878_));
 sky130_fd_sc_hd__a22oi_2 _19596_ (.A1(_11234_),
    .A2(_11275_),
    .B1(_11457_),
    .B2(\genblk1.pcpi_mul.rs1[12] ),
    .Y(_12879_));
 sky130_fd_sc_hd__or3_1 _19597_ (.A(_12877_),
    .B(_12878_),
    .C(_12879_),
    .X(_12880_));
 sky130_fd_sc_hd__o21ai_1 _19598_ (.A1(_12878_),
    .A2(_12879_),
    .B1(_12877_),
    .Y(_12881_));
 sky130_fd_sc_hd__o21bai_1 _19599_ (.A1(_12741_),
    .A2(_12743_),
    .B1_N(_12742_),
    .Y(_12882_));
 sky130_fd_sc_hd__and3_1 _19600_ (.A(_12880_),
    .B(_12881_),
    .C(_12882_),
    .X(_12883_));
 sky130_fd_sc_hd__a21o_1 _19601_ (.A1(_12880_),
    .A2(_12881_),
    .B1(_12882_),
    .X(_12884_));
 sky130_fd_sc_hd__and2b_1 _19602_ (.A_N(_12883_),
    .B(_12884_),
    .X(_12885_));
 sky130_fd_sc_hd__xnor2_1 _19603_ (.A(_12876_),
    .B(_12885_),
    .Y(_12886_));
 sky130_fd_sc_hd__nand2_1 _19604_ (.A(_12753_),
    .B(_12755_),
    .Y(_12887_));
 sky130_fd_sc_hd__a31o_1 _19605_ (.A1(_10805_),
    .A2(_11769_),
    .A3(_12783_),
    .B1(_12782_),
    .X(_12888_));
 sky130_fd_sc_hd__nand2_1 _19606_ (.A(_11066_),
    .B(\genblk1.pcpi_mul.rs2[15] ),
    .Y(_12889_));
 sky130_fd_sc_hd__nand4_2 _19607_ (.A(_10918_),
    .B(_11154_),
    .C(_11554_),
    .D(_11657_),
    .Y(_12890_));
 sky130_fd_sc_hd__a22o_1 _19608_ (.A1(\genblk1.pcpi_mul.rs1[10] ),
    .A2(_11661_),
    .B1(\genblk1.pcpi_mul.rs2[17] ),
    .B2(\genblk1.pcpi_mul.rs1[9] ),
    .X(_12891_));
 sky130_fd_sc_hd__nand3b_1 _19609_ (.A_N(_12889_),
    .B(_12890_),
    .C(_12891_),
    .Y(_12892_));
 sky130_fd_sc_hd__a21bo_1 _19610_ (.A1(_12890_),
    .A2(_12891_),
    .B1_N(_12889_),
    .X(_12893_));
 sky130_fd_sc_hd__nand3_1 _19611_ (.A(_12888_),
    .B(_12892_),
    .C(_12893_),
    .Y(_12894_));
 sky130_fd_sc_hd__a21o_1 _19612_ (.A1(_12892_),
    .A2(_12893_),
    .B1(_12888_),
    .X(_12895_));
 sky130_fd_sc_hd__nand3_1 _19613_ (.A(_12887_),
    .B(_12894_),
    .C(_12895_),
    .Y(_12896_));
 sky130_fd_sc_hd__a21o_1 _19614_ (.A1(_12894_),
    .A2(_12895_),
    .B1(_12887_),
    .X(_12897_));
 sky130_fd_sc_hd__a21bo_1 _19615_ (.A1(_12751_),
    .A2(_12758_),
    .B1_N(_12757_),
    .X(_12898_));
 sky130_fd_sc_hd__and3_1 _19616_ (.A(_12896_),
    .B(_12897_),
    .C(_12898_),
    .X(_12899_));
 sky130_fd_sc_hd__a21oi_1 _19617_ (.A1(_12896_),
    .A2(_12897_),
    .B1(_12898_),
    .Y(_12900_));
 sky130_fd_sc_hd__or3_4 _19618_ (.A(_12886_),
    .B(_12899_),
    .C(_12900_),
    .X(_12901_));
 sky130_fd_sc_hd__o21ai_1 _19619_ (.A1(_12899_),
    .A2(_12900_),
    .B1(_12886_),
    .Y(_12902_));
 sky130_fd_sc_hd__and3_1 _19620_ (.A(_12871_),
    .B(_12901_),
    .C(_12902_),
    .X(_12903_));
 sky130_fd_sc_hd__a21oi_1 _19621_ (.A1(_12901_),
    .A2(_12902_),
    .B1(_12871_),
    .Y(_12904_));
 sky130_fd_sc_hd__a211o_1 _19622_ (.A1(_12870_),
    .A2(_12764_),
    .B1(_12903_),
    .C1(_12904_),
    .X(_12905_));
 sky130_fd_sc_hd__o211ai_2 _19623_ (.A1(_12903_),
    .A2(_12904_),
    .B1(_12870_),
    .C1(_12764_),
    .Y(_12906_));
 sky130_fd_sc_hd__and2_1 _19624_ (.A(_12778_),
    .B(_12794_),
    .X(_12907_));
 sky130_fd_sc_hd__and4_1 _19625_ (.A(_10709_),
    .B(\genblk1.pcpi_mul.rs1[1] ),
    .C(\genblk1.pcpi_mul.rs2[25] ),
    .D(\genblk1.pcpi_mul.rs2[26] ),
    .X(_12908_));
 sky130_fd_sc_hd__clkbuf_2 _19626_ (.A(\genblk1.pcpi_mul.rs2[25] ),
    .X(_12909_));
 sky130_fd_sc_hd__clkbuf_2 _19627_ (.A(\genblk1.pcpi_mul.rs2[26] ),
    .X(_12910_));
 sky130_fd_sc_hd__a22oi_1 _19628_ (.A1(_10634_),
    .A2(_12909_),
    .B1(_12910_),
    .B2(_10709_),
    .Y(_12911_));
 sky130_fd_sc_hd__and4bb_1 _19629_ (.A_N(_12908_),
    .B_N(_12911_),
    .C(_10607_),
    .D(\genblk1.pcpi_mul.rs2[24] ),
    .X(_12912_));
 sky130_fd_sc_hd__o2bb2a_1 _19630_ (.A1_N(_11777_),
    .A2_N(\genblk1.pcpi_mul.rs2[24] ),
    .B1(_12908_),
    .B2(_12911_),
    .X(_12913_));
 sky130_fd_sc_hd__nor2_1 _19631_ (.A(_12912_),
    .B(_12913_),
    .Y(_12914_));
 sky130_fd_sc_hd__and2_1 _19632_ (.A(_12777_),
    .B(_12914_),
    .X(_12915_));
 sky130_fd_sc_hd__nor2_1 _19633_ (.A(_12777_),
    .B(_12914_),
    .Y(_12916_));
 sky130_fd_sc_hd__or2_1 _19634_ (.A(_12915_),
    .B(_12916_),
    .X(_12917_));
 sky130_fd_sc_hd__or2b_1 _19635_ (.A(_12791_),
    .B_N(_12790_),
    .X(_12918_));
 sky130_fd_sc_hd__nand2_1 _19636_ (.A(_12785_),
    .B(_12792_),
    .Y(_12919_));
 sky130_fd_sc_hd__nand2_1 _19637_ (.A(_11177_),
    .B(_11770_),
    .Y(_12920_));
 sky130_fd_sc_hd__and4_1 _19638_ (.A(_10756_),
    .B(\genblk1.pcpi_mul.rs1[7] ),
    .C(_12593_),
    .D(\genblk1.pcpi_mul.rs2[20] ),
    .X(_12921_));
 sky130_fd_sc_hd__a22o_1 _19639_ (.A1(_10851_),
    .A2(_12593_),
    .B1(_12232_),
    .B2(_10756_),
    .X(_12922_));
 sky130_fd_sc_hd__and2b_1 _19640_ (.A_N(_12921_),
    .B(_12922_),
    .X(_12923_));
 sky130_fd_sc_hd__xnor2_2 _19641_ (.A(_12920_),
    .B(_12923_),
    .Y(_12924_));
 sky130_fd_sc_hd__nand2_1 _19642_ (.A(_10794_),
    .B(\genblk1.pcpi_mul.rs2[21] ),
    .Y(_12925_));
 sky130_fd_sc_hd__and4_1 _19643_ (.A(\genblk1.pcpi_mul.rs1[3] ),
    .B(\genblk1.pcpi_mul.rs1[4] ),
    .C(\genblk1.pcpi_mul.rs2[22] ),
    .D(_12462_),
    .X(_12926_));
 sky130_fd_sc_hd__a22o_1 _19644_ (.A1(\genblk1.pcpi_mul.rs1[4] ),
    .A2(\genblk1.pcpi_mul.rs2[22] ),
    .B1(_12462_),
    .B2(\genblk1.pcpi_mul.rs1[3] ),
    .X(_12927_));
 sky130_fd_sc_hd__and2b_1 _19645_ (.A_N(_12926_),
    .B(_12927_),
    .X(_12928_));
 sky130_fd_sc_hd__xnor2_2 _19646_ (.A(_12925_),
    .B(_12928_),
    .Y(_12929_));
 sky130_fd_sc_hd__a31oi_4 _19647_ (.A1(_10721_),
    .A2(_12460_),
    .A3(_12788_),
    .B1(_12787_),
    .Y(_12930_));
 sky130_fd_sc_hd__xnor2_1 _19648_ (.A(_12929_),
    .B(_12930_),
    .Y(_12931_));
 sky130_fd_sc_hd__xnor2_1 _19649_ (.A(_12924_),
    .B(_12931_),
    .Y(_12932_));
 sky130_fd_sc_hd__a21oi_1 _19650_ (.A1(_12918_),
    .A2(_12919_),
    .B1(_12932_),
    .Y(_12933_));
 sky130_fd_sc_hd__and3_1 _19651_ (.A(_12918_),
    .B(_12919_),
    .C(_12932_),
    .X(_12934_));
 sky130_fd_sc_hd__or3_2 _19652_ (.A(_12917_),
    .B(_12933_),
    .C(_12934_),
    .X(_12935_));
 sky130_fd_sc_hd__o21ai_1 _19653_ (.A1(_12933_),
    .A2(_12934_),
    .B1(_12917_),
    .Y(_12936_));
 sky130_fd_sc_hd__nand3_1 _19654_ (.A(_12907_),
    .B(_12935_),
    .C(_12936_),
    .Y(_12937_));
 sky130_fd_sc_hd__a21o_1 _19655_ (.A1(_12935_),
    .A2(_12936_),
    .B1(_12907_),
    .X(_12938_));
 sky130_fd_sc_hd__and4_2 _19656_ (.A(_12905_),
    .B(_12906_),
    .C(_12937_),
    .D(_12938_),
    .X(_12939_));
 sky130_fd_sc_hd__a22oi_4 _19657_ (.A1(_12905_),
    .A2(_12906_),
    .B1(_12937_),
    .B2(_12938_),
    .Y(_12940_));
 sky130_fd_sc_hd__a211oi_2 _19658_ (.A1(_12869_),
    .A2(_12797_),
    .B1(_12939_),
    .C1(_12940_),
    .Y(_12941_));
 sky130_fd_sc_hd__o211a_1 _19659_ (.A1(_12939_),
    .A2(_12940_),
    .B1(_12869_),
    .C1(_12797_),
    .X(_12942_));
 sky130_fd_sc_hd__nor4_1 _19660_ (.A(_12867_),
    .B(_12868_),
    .C(_12941_),
    .D(_12942_),
    .Y(_12943_));
 sky130_fd_sc_hd__o22a_1 _19661_ (.A1(_12867_),
    .A2(_12868_),
    .B1(_12941_),
    .B2(_12942_),
    .X(_12944_));
 sky130_fd_sc_hd__a211oi_2 _19662_ (.A1(_12799_),
    .A2(_12801_),
    .B1(net345),
    .C1(_12944_),
    .Y(_12945_));
 sky130_fd_sc_hd__o211a_1 _19663_ (.A1(net346),
    .A2(_12944_),
    .B1(_12799_),
    .C1(_12801_),
    .X(_12946_));
 sky130_fd_sc_hd__or3_1 _19664_ (.A(_12820_),
    .B(_12945_),
    .C(_12946_),
    .X(_12947_));
 sky130_fd_sc_hd__o21ai_1 _19665_ (.A1(_12945_),
    .A2(_12946_),
    .B1(_12820_),
    .Y(_12948_));
 sky130_fd_sc_hd__o211a_1 _19666_ (.A1(_12803_),
    .A2(_12817_),
    .B1(_12947_),
    .C1(_12948_),
    .X(_12949_));
 sky130_fd_sc_hd__a211oi_1 _19667_ (.A1(_12947_),
    .A2(_12948_),
    .B1(_12803_),
    .C1(_12817_),
    .Y(_12950_));
 sky130_fd_sc_hd__or3_1 _19668_ (.A(_12679_),
    .B(_12949_),
    .C(_12950_),
    .X(_12951_));
 sky130_fd_sc_hd__o21ai_1 _19669_ (.A1(_12949_),
    .A2(_12950_),
    .B1(_12679_),
    .Y(_12952_));
 sky130_fd_sc_hd__o211a_1 _19670_ (.A1(_12807_),
    .A2(_12816_),
    .B1(_12951_),
    .C1(_12952_),
    .X(_12953_));
 sky130_fd_sc_hd__a211oi_2 _19671_ (.A1(_12951_),
    .A2(_12952_),
    .B1(_12807_),
    .C1(_12816_),
    .Y(_12954_));
 sky130_fd_sc_hd__nor2_1 _19672_ (.A(_12953_),
    .B(_12954_),
    .Y(_12955_));
 sky130_vsdinv _19673_ (.A(_12814_),
    .Y(_12956_));
 sky130_fd_sc_hd__and2b_1 _19674_ (.A_N(_12664_),
    .B(_12813_),
    .X(_12957_));
 sky130_fd_sc_hd__o32a_1 _19675_ (.A1(_12666_),
    .A2(_12674_),
    .A3(_12956_),
    .B1(_12957_),
    .B2(_12812_),
    .X(_12958_));
 sky130_fd_sc_hd__xnor2_1 _19676_ (.A(_12955_),
    .B(_12958_),
    .Y(_00072_));
 sky130_fd_sc_hd__a21o_1 _19677_ (.A1(_12731_),
    .A2(_12733_),
    .B1(_12819_),
    .X(_12959_));
 sky130_fd_sc_hd__nor3_1 _19678_ (.A(_12820_),
    .B(_12945_),
    .C(_12946_),
    .Y(_12960_));
 sky130_vsdinv _19679_ (.A(_12865_),
    .Y(_12961_));
 sky130_fd_sc_hd__nor2_1 _19680_ (.A(_12961_),
    .B(_12867_),
    .Y(_12962_));
 sky130_fd_sc_hd__nor2_1 _19681_ (.A(_12841_),
    .B(_12843_),
    .Y(_12963_));
 sky130_fd_sc_hd__xnor2_1 _19682_ (.A(_12962_),
    .B(_12963_),
    .Y(_12964_));
 sky130_vsdinv _19683_ (.A(_12941_),
    .Y(_12965_));
 sky130_fd_sc_hd__or4_1 _19684_ (.A(_12867_),
    .B(_12868_),
    .C(_12941_),
    .D(_12942_),
    .X(_12966_));
 sky130_fd_sc_hd__nand3_1 _19685_ (.A(_12871_),
    .B(_12901_),
    .C(_12902_),
    .Y(_12967_));
 sky130_fd_sc_hd__or2_1 _19686_ (.A(_12689_),
    .B(_12827_),
    .X(_12968_));
 sky130_fd_sc_hd__a211o_1 _19687_ (.A1(_12691_),
    .A2(_12826_),
    .B1(_12828_),
    .C1(_12831_),
    .X(_12969_));
 sky130_fd_sc_hd__or2b_1 _19688_ (.A(_12838_),
    .B_N(_12837_),
    .X(_12970_));
 sky130_fd_sc_hd__nand2_1 _19689_ (.A(_12832_),
    .B(_12839_),
    .Y(_12971_));
 sky130_fd_sc_hd__nand2_1 _19690_ (.A(_10639_),
    .B(\genblk1.pcpi_mul.rs1[26] ),
    .Y(_12972_));
 sky130_fd_sc_hd__clkbuf_4 _19691_ (.A(\genblk1.pcpi_mul.rs1[26] ),
    .X(_12973_));
 sky130_fd_sc_hd__nand2_1 _19692_ (.A(_10740_),
    .B(_12973_),
    .Y(_12974_));
 sky130_fd_sc_hd__nor2_1 _19693_ (.A(_12826_),
    .B(_12974_),
    .Y(_12975_));
 sky130_fd_sc_hd__a21oi_1 _19694_ (.A1(_12827_),
    .A2(_12972_),
    .B1(_12975_),
    .Y(_12976_));
 sky130_fd_sc_hd__buf_2 _19695_ (.A(_12546_),
    .X(_12977_));
 sky130_fd_sc_hd__nand2_2 _19696_ (.A(_10625_),
    .B(_12977_),
    .Y(_12978_));
 sky130_fd_sc_hd__xnor2_1 _19697_ (.A(_12976_),
    .B(_12978_),
    .Y(_12979_));
 sky130_fd_sc_hd__clkbuf_4 _19698_ (.A(\genblk1.pcpi_mul.rs1[27] ),
    .X(_12980_));
 sky130_fd_sc_hd__nand2_1 _19699_ (.A(_10695_),
    .B(_12980_),
    .Y(_12981_));
 sky130_fd_sc_hd__and4_1 _19700_ (.A(_10802_),
    .B(_10916_),
    .C(\genblk1.pcpi_mul.rs1[22] ),
    .D(\genblk1.pcpi_mul.rs1[23] ),
    .X(_12982_));
 sky130_fd_sc_hd__clkbuf_4 _19701_ (.A(\genblk1.pcpi_mul.rs1[22] ),
    .X(_12983_));
 sky130_fd_sc_hd__a22oi_2 _19702_ (.A1(_10702_),
    .A2(_12983_),
    .B1(_12537_),
    .B2(_11710_),
    .Y(_12984_));
 sky130_fd_sc_hd__nor2_1 _19703_ (.A(_12982_),
    .B(_12984_),
    .Y(_12985_));
 sky130_fd_sc_hd__xnor2_1 _19704_ (.A(_12981_),
    .B(_12985_),
    .Y(_12986_));
 sky130_fd_sc_hd__o21ba_1 _19705_ (.A1(_12833_),
    .A2(_12835_),
    .B1_N(_12834_),
    .X(_12987_));
 sky130_fd_sc_hd__xnor2_1 _19706_ (.A(_12986_),
    .B(_12987_),
    .Y(_12988_));
 sky130_fd_sc_hd__xnor2_1 _19707_ (.A(_12979_),
    .B(_12988_),
    .Y(_12989_));
 sky130_fd_sc_hd__a21oi_2 _19708_ (.A1(_12970_),
    .A2(_12971_),
    .B1(_12989_),
    .Y(_12990_));
 sky130_fd_sc_hd__and3_1 _19709_ (.A(_12970_),
    .B(_12971_),
    .C(_12989_),
    .X(_12991_));
 sky130_fd_sc_hd__a211oi_2 _19710_ (.A1(_12968_),
    .A2(_12969_),
    .B1(_12990_),
    .C1(_12991_),
    .Y(_12992_));
 sky130_fd_sc_hd__o211a_1 _19711_ (.A1(_12990_),
    .A2(_12991_),
    .B1(_12968_),
    .C1(_12969_),
    .X(_12993_));
 sky130_fd_sc_hd__nand3_2 _19712_ (.A(_12845_),
    .B(_12855_),
    .C(_12856_),
    .Y(_12994_));
 sky130_fd_sc_hd__a21o_1 _19713_ (.A1(_12876_),
    .A2(_12884_),
    .B1(_12883_),
    .X(_12995_));
 sky130_fd_sc_hd__nand2_1 _19714_ (.A(_12849_),
    .B(_12851_),
    .Y(_12996_));
 sky130_fd_sc_hd__a31o_1 _19715_ (.A1(_10960_),
    .A2(_12285_),
    .A3(_12874_),
    .B1(_12873_),
    .X(_12997_));
 sky130_fd_sc_hd__nand4_2 _19716_ (.A(_10997_),
    .B(_11085_),
    .C(_12069_),
    .D(_12078_),
    .Y(_12998_));
 sky130_fd_sc_hd__a22o_1 _19717_ (.A1(_11195_),
    .A2(_11957_),
    .B1(_12143_),
    .B2(_10995_),
    .X(_12999_));
 sky130_fd_sc_hd__nand4_2 _19718_ (.A(_10736_),
    .B(_12154_),
    .C(_12998_),
    .D(_12999_),
    .Y(_13000_));
 sky130_fd_sc_hd__a22o_1 _19719_ (.A1(_10993_),
    .A2(_12271_),
    .B1(_12998_),
    .B2(_12999_),
    .X(_13001_));
 sky130_fd_sc_hd__nand3_2 _19720_ (.A(_12997_),
    .B(_13000_),
    .C(_13001_),
    .Y(_13002_));
 sky130_fd_sc_hd__a21o_1 _19721_ (.A1(_13000_),
    .A2(_13001_),
    .B1(_12997_),
    .X(_13003_));
 sky130_fd_sc_hd__nand3_2 _19722_ (.A(_12996_),
    .B(_13002_),
    .C(_13003_),
    .Y(_13004_));
 sky130_fd_sc_hd__a21o_1 _19723_ (.A1(_13002_),
    .A2(_13003_),
    .B1(_12996_),
    .X(_13005_));
 sky130_fd_sc_hd__and3_2 _19724_ (.A(_12995_),
    .B(_13004_),
    .C(_13005_),
    .X(_13006_));
 sky130_fd_sc_hd__a21oi_2 _19725_ (.A1(_13004_),
    .A2(_13005_),
    .B1(_12995_),
    .Y(_13007_));
 sky130_fd_sc_hd__a211oi_4 _19726_ (.A1(_12853_),
    .A2(_12855_),
    .B1(_13006_),
    .C1(_13007_),
    .Y(_13008_));
 sky130_fd_sc_hd__o211a_1 _19727_ (.A1(_13006_),
    .A2(_13007_),
    .B1(_12853_),
    .C1(_12855_),
    .X(_13009_));
 sky130_fd_sc_hd__a211oi_4 _19728_ (.A1(_12994_),
    .A2(_12859_),
    .B1(_13008_),
    .C1(_13009_),
    .Y(_13010_));
 sky130_fd_sc_hd__o211a_1 _19729_ (.A1(_13008_),
    .A2(_13009_),
    .B1(_12994_),
    .C1(_12859_),
    .X(_13011_));
 sky130_fd_sc_hd__nor4_1 _19730_ (.A(_12992_),
    .B(_12993_),
    .C(_13010_),
    .D(_13011_),
    .Y(_13012_));
 sky130_fd_sc_hd__o22a_1 _19731_ (.A1(_12992_),
    .A2(_12993_),
    .B1(_13010_),
    .B2(_13011_),
    .X(_13013_));
 sky130_fd_sc_hd__a211oi_1 _19732_ (.A1(_12967_),
    .A2(_12905_),
    .B1(net419),
    .C1(_13013_),
    .Y(_13014_));
 sky130_fd_sc_hd__o211a_1 _19733_ (.A1(net419),
    .A2(_13013_),
    .B1(_12967_),
    .C1(_12905_),
    .X(_13015_));
 sky130_fd_sc_hd__a211oi_1 _19734_ (.A1(_12861_),
    .A2(_12863_),
    .B1(_13014_),
    .C1(_13015_),
    .Y(_13016_));
 sky130_fd_sc_hd__o211a_1 _19735_ (.A1(_13014_),
    .A2(_13015_),
    .B1(_12861_),
    .C1(_12863_),
    .X(_13017_));
 sky130_fd_sc_hd__and3_1 _19736_ (.A(_12907_),
    .B(_12935_),
    .C(_12936_),
    .X(_13018_));
 sky130_fd_sc_hd__nand3_2 _19737_ (.A(_12896_),
    .B(_12897_),
    .C(_12898_),
    .Y(_13019_));
 sky130_fd_sc_hd__nand2_1 _19738_ (.A(_10960_),
    .B(_11830_),
    .Y(_13020_));
 sky130_fd_sc_hd__and4_1 _19739_ (.A(_11140_),
    .B(_11143_),
    .C(_11697_),
    .D(_12714_),
    .X(_13021_));
 sky130_fd_sc_hd__a22o_1 _19740_ (.A1(_11106_),
    .A2(_11697_),
    .B1(_12714_),
    .B2(_11140_),
    .X(_13022_));
 sky130_fd_sc_hd__and2b_1 _19741_ (.A_N(_13021_),
    .B(_13022_),
    .X(_13023_));
 sky130_fd_sc_hd__xnor2_1 _19742_ (.A(_13020_),
    .B(_13023_),
    .Y(_13024_));
 sky130_fd_sc_hd__nand2_1 _19743_ (.A(\genblk1.pcpi_mul.rs2[12] ),
    .B(_11588_),
    .Y(_13025_));
 sky130_fd_sc_hd__and4_1 _19744_ (.A(_11239_),
    .B(\genblk1.pcpi_mul.rs1[13] ),
    .C(_11352_),
    .D(\genblk1.pcpi_mul.rs1[14] ),
    .X(_13026_));
 sky130_fd_sc_hd__a22oi_2 _19745_ (.A1(_11275_),
    .A2(_11457_),
    .B1(_11480_),
    .B2(_11239_),
    .Y(_13027_));
 sky130_fd_sc_hd__or3_1 _19746_ (.A(_13025_),
    .B(_13026_),
    .C(_13027_),
    .X(_13028_));
 sky130_fd_sc_hd__o21ai_1 _19747_ (.A1(_13026_),
    .A2(_13027_),
    .B1(_13025_),
    .Y(_13029_));
 sky130_fd_sc_hd__o21bai_1 _19748_ (.A1(_12877_),
    .A2(_12879_),
    .B1_N(_12878_),
    .Y(_13030_));
 sky130_fd_sc_hd__and3_1 _19749_ (.A(_13028_),
    .B(_13029_),
    .C(_13030_),
    .X(_13031_));
 sky130_fd_sc_hd__a21o_1 _19750_ (.A1(_13028_),
    .A2(_13029_),
    .B1(_13030_),
    .X(_13032_));
 sky130_fd_sc_hd__and2b_1 _19751_ (.A_N(_13031_),
    .B(_13032_),
    .X(_13033_));
 sky130_fd_sc_hd__xnor2_1 _19752_ (.A(_13024_),
    .B(_13033_),
    .Y(_13034_));
 sky130_fd_sc_hd__nand2_1 _19753_ (.A(_12890_),
    .B(_12892_),
    .Y(_13035_));
 sky130_fd_sc_hd__a31o_1 _19754_ (.A1(_10858_),
    .A2(_11769_),
    .A3(_12922_),
    .B1(_12921_),
    .X(_13036_));
 sky130_fd_sc_hd__nand4_2 _19755_ (.A(_11154_),
    .B(_11066_),
    .C(_11661_),
    .D(_11657_),
    .Y(_13037_));
 sky130_fd_sc_hd__a22o_1 _19756_ (.A1(\genblk1.pcpi_mul.rs1[11] ),
    .A2(_11661_),
    .B1(\genblk1.pcpi_mul.rs2[17] ),
    .B2(\genblk1.pcpi_mul.rs1[10] ),
    .X(_13038_));
 sky130_fd_sc_hd__nand4_1 _19757_ (.A(_11260_),
    .B(_12364_),
    .C(_13037_),
    .D(_13038_),
    .Y(_13039_));
 sky130_fd_sc_hd__a22o_1 _19758_ (.A1(_12098_),
    .A2(_12364_),
    .B1(_13037_),
    .B2(_13038_),
    .X(_13040_));
 sky130_fd_sc_hd__nand3_1 _19759_ (.A(_13036_),
    .B(_13039_),
    .C(_13040_),
    .Y(_13041_));
 sky130_fd_sc_hd__a21o_1 _19760_ (.A1(_13039_),
    .A2(_13040_),
    .B1(_13036_),
    .X(_13042_));
 sky130_fd_sc_hd__nand3_1 _19761_ (.A(_13035_),
    .B(_13041_),
    .C(_13042_),
    .Y(_13043_));
 sky130_fd_sc_hd__a21o_1 _19762_ (.A1(_13041_),
    .A2(_13042_),
    .B1(_13035_),
    .X(_13044_));
 sky130_fd_sc_hd__a21bo_1 _19763_ (.A1(_12887_),
    .A2(_12895_),
    .B1_N(_12894_),
    .X(_13045_));
 sky130_fd_sc_hd__and3_1 _19764_ (.A(_13043_),
    .B(_13044_),
    .C(_13045_),
    .X(_13046_));
 sky130_fd_sc_hd__a21oi_1 _19765_ (.A1(_13043_),
    .A2(_13044_),
    .B1(_13045_),
    .Y(_13047_));
 sky130_fd_sc_hd__or3_2 _19766_ (.A(_13034_),
    .B(_13046_),
    .C(_13047_),
    .X(_13048_));
 sky130_fd_sc_hd__o21ai_1 _19767_ (.A1(_13046_),
    .A2(_13047_),
    .B1(_13034_),
    .Y(_13049_));
 sky130_fd_sc_hd__and3_2 _19768_ (.A(_12933_),
    .B(_13048_),
    .C(_13049_),
    .X(_13050_));
 sky130_fd_sc_hd__a21oi_2 _19769_ (.A1(_13048_),
    .A2(_13049_),
    .B1(_12933_),
    .Y(_13051_));
 sky130_fd_sc_hd__a211oi_4 _19770_ (.A1(_13019_),
    .A2(_12901_),
    .B1(_13050_),
    .C1(_13051_),
    .Y(_13052_));
 sky130_fd_sc_hd__o211a_1 _19771_ (.A1(_13050_),
    .A2(_13051_),
    .B1(_13019_),
    .C1(_12901_),
    .X(_13053_));
 sky130_fd_sc_hd__clkbuf_2 _19772_ (.A(\genblk1.pcpi_mul.rs2[27] ),
    .X(_13054_));
 sky130_fd_sc_hd__clkbuf_2 _19773_ (.A(_13054_),
    .X(_13055_));
 sky130_fd_sc_hd__clkbuf_4 _19774_ (.A(_13055_),
    .X(_13056_));
 sky130_fd_sc_hd__nand2_2 _19775_ (.A(_10623_),
    .B(_13056_),
    .Y(_13057_));
 sky130_fd_sc_hd__nand2_1 _19776_ (.A(_10649_),
    .B(_12775_),
    .Y(_13058_));
 sky130_fd_sc_hd__and4_1 _19777_ (.A(_10634_),
    .B(_10628_),
    .C(_12770_),
    .D(_12910_),
    .X(_13059_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19778_ (.A(_12909_),
    .X(_13060_));
 sky130_fd_sc_hd__clkbuf_2 _19779_ (.A(\genblk1.pcpi_mul.rs2[26] ),
    .X(_13061_));
 sky130_fd_sc_hd__a22oi_2 _19780_ (.A1(_10607_),
    .A2(_13060_),
    .B1(_13061_),
    .B2(_10786_),
    .Y(_13062_));
 sky130_fd_sc_hd__nor2_1 _19781_ (.A(_13059_),
    .B(_13062_),
    .Y(_13063_));
 sky130_fd_sc_hd__xnor2_1 _19782_ (.A(_13058_),
    .B(_13063_),
    .Y(_13064_));
 sky130_fd_sc_hd__nor2_1 _19783_ (.A(_12908_),
    .B(_12912_),
    .Y(_13065_));
 sky130_fd_sc_hd__xnor2_1 _19784_ (.A(_13064_),
    .B(_13065_),
    .Y(_13066_));
 sky130_fd_sc_hd__xnor2_1 _19785_ (.A(_13057_),
    .B(_13066_),
    .Y(_13067_));
 sky130_fd_sc_hd__and2b_1 _19786_ (.A_N(_12930_),
    .B(_12929_),
    .X(_13068_));
 sky130_fd_sc_hd__a21o_1 _19787_ (.A1(_12924_),
    .A2(_12931_),
    .B1(_13068_),
    .X(_13069_));
 sky130_fd_sc_hd__nand2_1 _19788_ (.A(_11280_),
    .B(_11894_),
    .Y(_13070_));
 sky130_fd_sc_hd__and4_1 _19789_ (.A(_10851_),
    .B(_10907_),
    .C(_12333_),
    .D(_12232_),
    .X(_13071_));
 sky130_fd_sc_hd__a22o_1 _19790_ (.A1(_10907_),
    .A2(_12333_),
    .B1(_12020_),
    .B2(_10851_),
    .X(_13072_));
 sky130_fd_sc_hd__and2b_1 _19791_ (.A_N(_13071_),
    .B(_13072_),
    .X(_13073_));
 sky130_fd_sc_hd__xnor2_1 _19792_ (.A(_13070_),
    .B(_13073_),
    .Y(_13074_));
 sky130_fd_sc_hd__and2_1 _19793_ (.A(_10978_),
    .B(\genblk1.pcpi_mul.rs2[21] ),
    .X(_13075_));
 sky130_fd_sc_hd__nand4_2 _19794_ (.A(_10741_),
    .B(_10745_),
    .C(_12327_),
    .D(_12464_),
    .Y(_13076_));
 sky130_fd_sc_hd__a22o_1 _19795_ (.A1(_10793_),
    .A2(_12321_),
    .B1(_12464_),
    .B2(_10718_),
    .X(_13077_));
 sky130_fd_sc_hd__nand3_1 _19796_ (.A(_13075_),
    .B(_13076_),
    .C(_13077_),
    .Y(_13078_));
 sky130_fd_sc_hd__a21o_1 _19797_ (.A1(_13076_),
    .A2(_13077_),
    .B1(_13075_),
    .X(_13079_));
 sky130_fd_sc_hd__a31o_1 _19798_ (.A1(_10790_),
    .A2(_12460_),
    .A3(_12927_),
    .B1(_12926_),
    .X(_13080_));
 sky130_fd_sc_hd__nand3_1 _19799_ (.A(_13078_),
    .B(_13079_),
    .C(_13080_),
    .Y(_13081_));
 sky130_fd_sc_hd__a21o_1 _19800_ (.A1(_13078_),
    .A2(_13079_),
    .B1(_13080_),
    .X(_13082_));
 sky130_fd_sc_hd__nand3_1 _19801_ (.A(_13074_),
    .B(_13081_),
    .C(_13082_),
    .Y(_13083_));
 sky130_fd_sc_hd__a21o_1 _19802_ (.A1(_13081_),
    .A2(_13082_),
    .B1(_13074_),
    .X(_13084_));
 sky130_fd_sc_hd__nand3_2 _19803_ (.A(_12915_),
    .B(_13083_),
    .C(_13084_),
    .Y(_13085_));
 sky130_fd_sc_hd__a21o_1 _19804_ (.A1(_13083_),
    .A2(_13084_),
    .B1(_12915_),
    .X(_13086_));
 sky130_fd_sc_hd__nand3_2 _19805_ (.A(_13069_),
    .B(_13085_),
    .C(_13086_),
    .Y(_13087_));
 sky130_fd_sc_hd__a21o_1 _19806_ (.A1(_13085_),
    .A2(_13086_),
    .B1(_13069_),
    .X(_13088_));
 sky130_fd_sc_hd__and3_1 _19807_ (.A(_13067_),
    .B(_13087_),
    .C(_13088_),
    .X(_13089_));
 sky130_fd_sc_hd__a21oi_1 _19808_ (.A1(_13087_),
    .A2(_13088_),
    .B1(_13067_),
    .Y(_13090_));
 sky130_fd_sc_hd__or3_1 _19809_ (.A(_12935_),
    .B(_13089_),
    .C(_13090_),
    .X(_13091_));
 sky130_fd_sc_hd__o21ai_1 _19810_ (.A1(_13089_),
    .A2(_13090_),
    .B1(_12935_),
    .Y(_13092_));
 sky130_fd_sc_hd__or4bb_2 _19811_ (.A(_13052_),
    .B(_13053_),
    .C_N(_13091_),
    .D_N(_13092_),
    .X(_13093_));
 sky130_fd_sc_hd__a2bb2o_1 _19812_ (.A1_N(_13052_),
    .A2_N(_13053_),
    .B1(_13091_),
    .B2(_13092_),
    .X(_13094_));
 sky130_fd_sc_hd__o211a_1 _19813_ (.A1(_13018_),
    .A2(_12939_),
    .B1(_13093_),
    .C1(_13094_),
    .X(_13095_));
 sky130_fd_sc_hd__a211oi_1 _19814_ (.A1(_13093_),
    .A2(_13094_),
    .B1(_13018_),
    .C1(_12939_),
    .Y(_13096_));
 sky130_fd_sc_hd__nor4_1 _19815_ (.A(_13016_),
    .B(_13017_),
    .C(_13095_),
    .D(_13096_),
    .Y(_13097_));
 sky130_fd_sc_hd__o22a_1 _19816_ (.A1(_13016_),
    .A2(_13017_),
    .B1(_13095_),
    .B2(_13096_),
    .X(_13098_));
 sky130_fd_sc_hd__a211oi_2 _19817_ (.A1(_12965_),
    .A2(_12966_),
    .B1(net344),
    .C1(_13098_),
    .Y(_13099_));
 sky130_fd_sc_hd__o211a_1 _19818_ (.A1(net344),
    .A2(_13098_),
    .B1(_12965_),
    .C1(_12966_),
    .X(_13100_));
 sky130_fd_sc_hd__or3_1 _19819_ (.A(_12964_),
    .B(_13099_),
    .C(_13100_),
    .X(_13101_));
 sky130_fd_sc_hd__o21ai_1 _19820_ (.A1(_13099_),
    .A2(_13100_),
    .B1(_12964_),
    .Y(_13102_));
 sky130_fd_sc_hd__o211a_1 _19821_ (.A1(_12945_),
    .A2(_12960_),
    .B1(_13101_),
    .C1(_13102_),
    .X(_13103_));
 sky130_fd_sc_hd__a211oi_1 _19822_ (.A1(_13101_),
    .A2(_13102_),
    .B1(_12945_),
    .C1(_12960_),
    .Y(_13104_));
 sky130_fd_sc_hd__or3_1 _19823_ (.A(_12959_),
    .B(_13103_),
    .C(_13104_),
    .X(_13105_));
 sky130_fd_sc_hd__o21ai_1 _19824_ (.A1(_13103_),
    .A2(_13104_),
    .B1(_12959_),
    .Y(_13106_));
 sky130_fd_sc_hd__nor3_1 _19825_ (.A(_12679_),
    .B(_12949_),
    .C(_12950_),
    .Y(_13107_));
 sky130_fd_sc_hd__a211oi_1 _19826_ (.A1(_13105_),
    .A2(_13106_),
    .B1(_12949_),
    .C1(_13107_),
    .Y(_13108_));
 sky130_fd_sc_hd__o211a_1 _19827_ (.A1(_12949_),
    .A2(_13107_),
    .B1(_13105_),
    .C1(_13106_),
    .X(_13109_));
 sky130_fd_sc_hd__nor2_1 _19828_ (.A(_13108_),
    .B(_13109_),
    .Y(_13110_));
 sky130_fd_sc_hd__o21ba_1 _19829_ (.A1(_12954_),
    .A2(_12958_),
    .B1_N(_12953_),
    .X(_13111_));
 sky130_fd_sc_hd__xnor2_1 _19830_ (.A(_13110_),
    .B(_13111_),
    .Y(_00073_));
 sky130_fd_sc_hd__or2_1 _19831_ (.A(_12962_),
    .B(_12963_),
    .X(_13112_));
 sky130_fd_sc_hd__nor3_1 _19832_ (.A(_12964_),
    .B(_13099_),
    .C(_13100_),
    .Y(_13113_));
 sky130_fd_sc_hd__or2_1 _19833_ (.A(_13014_),
    .B(_13016_),
    .X(_13114_));
 sky130_fd_sc_hd__nor2_1 _19834_ (.A(_12990_),
    .B(_12992_),
    .Y(_13115_));
 sky130_fd_sc_hd__xor2_1 _19835_ (.A(_13114_),
    .B(_13115_),
    .X(_13116_));
 sky130_fd_sc_hd__or2_1 _19836_ (.A(_12826_),
    .B(_12974_),
    .X(_13117_));
 sky130_fd_sc_hd__a211o_1 _19837_ (.A1(_12827_),
    .A2(_12972_),
    .B1(_12978_),
    .C1(_12975_),
    .X(_13118_));
 sky130_fd_sc_hd__or2b_1 _19838_ (.A(_12987_),
    .B_N(_12986_),
    .X(_13119_));
 sky130_fd_sc_hd__nand2_1 _19839_ (.A(_12979_),
    .B(_12988_),
    .Y(_13120_));
 sky130_fd_sc_hd__nand2_1 _19840_ (.A(_10747_),
    .B(_12980_),
    .Y(_13121_));
 sky130_fd_sc_hd__nand2_2 _19841_ (.A(_10610_),
    .B(\genblk1.pcpi_mul.rs1[27] ),
    .Y(_13122_));
 sky130_fd_sc_hd__nor2_1 _19842_ (.A(_12972_),
    .B(_13122_),
    .Y(_13123_));
 sky130_fd_sc_hd__a21oi_1 _19843_ (.A1(_12974_),
    .A2(_13121_),
    .B1(_13123_),
    .Y(_13124_));
 sky130_fd_sc_hd__buf_2 _19844_ (.A(_12700_),
    .X(_13125_));
 sky130_fd_sc_hd__nand2_2 _19845_ (.A(_10644_),
    .B(_13125_),
    .Y(_13126_));
 sky130_fd_sc_hd__xnor2_1 _19846_ (.A(_13124_),
    .B(_13126_),
    .Y(_13127_));
 sky130_fd_sc_hd__clkbuf_4 _19847_ (.A(\genblk1.pcpi_mul.rs1[28] ),
    .X(_13128_));
 sky130_fd_sc_hd__nand2_1 _19848_ (.A(_10695_),
    .B(_13128_),
    .Y(_13129_));
 sky130_fd_sc_hd__and4_1 _19849_ (.A(_10699_),
    .B(_10706_),
    .C(\genblk1.pcpi_mul.rs1[23] ),
    .D(\genblk1.pcpi_mul.rs1[24] ),
    .X(_13130_));
 sky130_fd_sc_hd__a22oi_2 _19850_ (.A1(_10707_),
    .A2(\genblk1.pcpi_mul.rs1[23] ),
    .B1(\genblk1.pcpi_mul.rs1[24] ),
    .B2(_10802_),
    .Y(_13131_));
 sky130_fd_sc_hd__nor2_1 _19851_ (.A(_13130_),
    .B(_13131_),
    .Y(_13132_));
 sky130_fd_sc_hd__xnor2_2 _19852_ (.A(_13129_),
    .B(_13132_),
    .Y(_13133_));
 sky130_fd_sc_hd__o21ba_1 _19853_ (.A1(_12981_),
    .A2(_12984_),
    .B1_N(_12982_),
    .X(_13134_));
 sky130_fd_sc_hd__xnor2_1 _19854_ (.A(_13133_),
    .B(_13134_),
    .Y(_13135_));
 sky130_fd_sc_hd__xnor2_1 _19855_ (.A(_13127_),
    .B(_13135_),
    .Y(_13136_));
 sky130_fd_sc_hd__a21oi_1 _19856_ (.A1(_13119_),
    .A2(_13120_),
    .B1(_13136_),
    .Y(_13137_));
 sky130_fd_sc_hd__and3_1 _19857_ (.A(_13119_),
    .B(_13120_),
    .C(_13136_),
    .X(_13138_));
 sky130_fd_sc_hd__a211oi_1 _19858_ (.A1(_13117_),
    .A2(_13118_),
    .B1(_13137_),
    .C1(_13138_),
    .Y(_13139_));
 sky130_fd_sc_hd__o211a_1 _19859_ (.A1(_13137_),
    .A2(_13138_),
    .B1(_13117_),
    .C1(_13118_),
    .X(_13140_));
 sky130_fd_sc_hd__a21o_1 _19860_ (.A1(_13024_),
    .A2(_13032_),
    .B1(_13031_),
    .X(_13141_));
 sky130_fd_sc_hd__nand2_1 _19861_ (.A(_12998_),
    .B(_13000_),
    .Y(_13142_));
 sky130_fd_sc_hd__a31o_1 _19862_ (.A1(_11189_),
    .A2(_11946_),
    .A3(_13022_),
    .B1(_13021_),
    .X(_13143_));
 sky130_fd_sc_hd__nand2_1 _19863_ (.A(_10735_),
    .B(_12281_),
    .Y(_13144_));
 sky130_fd_sc_hd__nand4_2 _19864_ (.A(_12172_),
    .B(_10837_),
    .C(_12143_),
    .D(_12153_),
    .Y(_13145_));
 sky130_fd_sc_hd__a22o_1 _19865_ (.A1(_10839_),
    .A2(_12143_),
    .B1(_12153_),
    .B2(_10836_),
    .X(_13146_));
 sky130_fd_sc_hd__nand3b_1 _19866_ (.A_N(_13144_),
    .B(_13145_),
    .C(_13146_),
    .Y(_13147_));
 sky130_fd_sc_hd__a21bo_1 _19867_ (.A1(_13145_),
    .A2(_13146_),
    .B1_N(_13144_),
    .X(_13148_));
 sky130_fd_sc_hd__nand3_2 _19868_ (.A(_13143_),
    .B(_13147_),
    .C(_13148_),
    .Y(_13149_));
 sky130_fd_sc_hd__a21o_1 _19869_ (.A1(_13147_),
    .A2(_13148_),
    .B1(_13143_),
    .X(_13150_));
 sky130_fd_sc_hd__nand3_2 _19870_ (.A(_13142_),
    .B(_13149_),
    .C(_13150_),
    .Y(_13151_));
 sky130_fd_sc_hd__a21o_1 _19871_ (.A1(_13149_),
    .A2(_13150_),
    .B1(_13142_),
    .X(_13152_));
 sky130_fd_sc_hd__and3_1 _19872_ (.A(_13141_),
    .B(_13151_),
    .C(_13152_),
    .X(_13153_));
 sky130_fd_sc_hd__a21oi_1 _19873_ (.A1(_13151_),
    .A2(_13152_),
    .B1(_13141_),
    .Y(_13154_));
 sky130_fd_sc_hd__a211o_2 _19874_ (.A1(_13002_),
    .A2(_13004_),
    .B1(_13153_),
    .C1(_13154_),
    .X(_13155_));
 sky130_fd_sc_hd__o211ai_2 _19875_ (.A1(_13153_),
    .A2(_13154_),
    .B1(_13002_),
    .C1(_13004_),
    .Y(_13156_));
 sky130_fd_sc_hd__o211ai_2 _19876_ (.A1(_13006_),
    .A2(_13008_),
    .B1(_13155_),
    .C1(_13156_),
    .Y(_13157_));
 sky130_fd_sc_hd__a211o_1 _19877_ (.A1(_13155_),
    .A2(_13156_),
    .B1(_13006_),
    .C1(_13008_),
    .X(_13158_));
 sky130_fd_sc_hd__or4bb_2 _19878_ (.A(_13139_),
    .B(_13140_),
    .C_N(_13157_),
    .D_N(_13158_),
    .X(_13159_));
 sky130_fd_sc_hd__a2bb2o_1 _19879_ (.A1_N(_13139_),
    .A2_N(_13140_),
    .B1(_13157_),
    .B2(_13158_),
    .X(_13160_));
 sky130_fd_sc_hd__o211ai_4 _19880_ (.A1(_13050_),
    .A2(_13052_),
    .B1(_13159_),
    .C1(_13160_),
    .Y(_13161_));
 sky130_fd_sc_hd__a211o_1 _19881_ (.A1(_13159_),
    .A2(_13160_),
    .B1(_13050_),
    .C1(_13052_),
    .X(_13162_));
 sky130_fd_sc_hd__o211ai_4 _19882_ (.A1(_13010_),
    .A2(net363),
    .B1(_13161_),
    .C1(_13162_),
    .Y(_13163_));
 sky130_fd_sc_hd__a211o_1 _19883_ (.A1(_13161_),
    .A2(_13162_),
    .B1(_13010_),
    .C1(net364),
    .X(_13164_));
 sky130_fd_sc_hd__nand3_1 _19884_ (.A(_13043_),
    .B(_13044_),
    .C(_13045_),
    .Y(_13165_));
 sky130_fd_sc_hd__nand2_1 _19885_ (.A(_11900_),
    .B(_12070_),
    .Y(_13166_));
 sky130_fd_sc_hd__and4_1 _19886_ (.A(_10962_),
    .B(_11106_),
    .C(_12714_),
    .D(_11829_),
    .X(_13167_));
 sky130_fd_sc_hd__a22o_1 _19887_ (.A1(_11905_),
    .A2(_12714_),
    .B1(_11829_),
    .B2(_10962_),
    .X(_13168_));
 sky130_fd_sc_hd__and2b_1 _19888_ (.A_N(_13167_),
    .B(_13168_),
    .X(_13169_));
 sky130_fd_sc_hd__xnor2_2 _19889_ (.A(_13166_),
    .B(_13169_),
    .Y(_13170_));
 sky130_fd_sc_hd__nand2_1 _19890_ (.A(_11349_),
    .B(_11597_),
    .Y(_13171_));
 sky130_fd_sc_hd__and4_1 _19891_ (.A(_11240_),
    .B(_11910_),
    .C(_11480_),
    .D(_11588_),
    .X(_13172_));
 sky130_fd_sc_hd__a22oi_2 _19892_ (.A1(_11353_),
    .A2(_11379_),
    .B1(_11488_),
    .B2(_11795_),
    .Y(_13173_));
 sky130_fd_sc_hd__or3_1 _19893_ (.A(_13171_),
    .B(_13172_),
    .C(_13173_),
    .X(_13174_));
 sky130_fd_sc_hd__o21ai_1 _19894_ (.A1(_13172_),
    .A2(_13173_),
    .B1(_13171_),
    .Y(_13175_));
 sky130_fd_sc_hd__o21bai_2 _19895_ (.A1(_13025_),
    .A2(_13027_),
    .B1_N(_13026_),
    .Y(_13176_));
 sky130_fd_sc_hd__and3_1 _19896_ (.A(_13174_),
    .B(_13175_),
    .C(_13176_),
    .X(_13177_));
 sky130_fd_sc_hd__a21o_1 _19897_ (.A1(_13174_),
    .A2(_13175_),
    .B1(_13176_),
    .X(_13178_));
 sky130_fd_sc_hd__and2b_1 _19898_ (.A_N(_13177_),
    .B(_13178_),
    .X(_13179_));
 sky130_fd_sc_hd__xnor2_1 _19899_ (.A(_13170_),
    .B(_13179_),
    .Y(_13180_));
 sky130_fd_sc_hd__nand2_1 _19900_ (.A(_13037_),
    .B(_13039_),
    .Y(_13181_));
 sky130_fd_sc_hd__a31o_1 _19901_ (.A1(_11036_),
    .A2(_11894_),
    .A3(_13072_),
    .B1(_13071_),
    .X(_13182_));
 sky130_fd_sc_hd__nand2_1 _19902_ (.A(_11712_),
    .B(_12364_),
    .Y(_13183_));
 sky130_fd_sc_hd__nand4_2 _19903_ (.A(_11054_),
    .B(_12098_),
    .C(_11922_),
    .D(_11780_),
    .Y(_13184_));
 sky130_fd_sc_hd__a22o_1 _19904_ (.A1(_11170_),
    .A2(_11922_),
    .B1(_11780_),
    .B2(_11066_),
    .X(_13185_));
 sky130_fd_sc_hd__nand3b_1 _19905_ (.A_N(_13183_),
    .B(_13184_),
    .C(_13185_),
    .Y(_13186_));
 sky130_fd_sc_hd__a21bo_1 _19906_ (.A1(_13184_),
    .A2(_13185_),
    .B1_N(_13183_),
    .X(_13187_));
 sky130_fd_sc_hd__nand3_1 _19907_ (.A(_13182_),
    .B(_13186_),
    .C(_13187_),
    .Y(_13188_));
 sky130_fd_sc_hd__a21o_1 _19908_ (.A1(_13186_),
    .A2(_13187_),
    .B1(_13182_),
    .X(_13189_));
 sky130_fd_sc_hd__nand3_1 _19909_ (.A(_13181_),
    .B(_13188_),
    .C(_13189_),
    .Y(_13190_));
 sky130_fd_sc_hd__a21o_1 _19910_ (.A1(_13188_),
    .A2(_13189_),
    .B1(_13181_),
    .X(_13191_));
 sky130_fd_sc_hd__a21bo_1 _19911_ (.A1(_13035_),
    .A2(_13042_),
    .B1_N(_13041_),
    .X(_13192_));
 sky130_fd_sc_hd__and3_1 _19912_ (.A(_13190_),
    .B(_13191_),
    .C(_13192_),
    .X(_13193_));
 sky130_fd_sc_hd__a21oi_1 _19913_ (.A1(_13190_),
    .A2(_13191_),
    .B1(_13192_),
    .Y(_13194_));
 sky130_fd_sc_hd__nor3_1 _19914_ (.A(_13180_),
    .B(_13193_),
    .C(_13194_),
    .Y(_13195_));
 sky130_fd_sc_hd__o21a_1 _19915_ (.A1(_13193_),
    .A2(_13194_),
    .B1(_13180_),
    .X(_13196_));
 sky130_fd_sc_hd__a211oi_1 _19916_ (.A1(_13085_),
    .A2(_13087_),
    .B1(net366),
    .C1(_13196_),
    .Y(_13197_));
 sky130_fd_sc_hd__o211a_1 _19917_ (.A1(net366),
    .A2(_13196_),
    .B1(_13085_),
    .C1(_13087_),
    .X(_13198_));
 sky130_fd_sc_hd__a211o_1 _19918_ (.A1(_13165_),
    .A2(_13048_),
    .B1(_13197_),
    .C1(_13198_),
    .X(_13199_));
 sky130_fd_sc_hd__o211ai_2 _19919_ (.A1(_13197_),
    .A2(_13198_),
    .B1(_13165_),
    .C1(_13048_),
    .Y(_13200_));
 sky130_fd_sc_hd__nand2_1 _19920_ (.A(_13081_),
    .B(_13083_),
    .Y(_13201_));
 sky130_fd_sc_hd__and2b_1 _19921_ (.A_N(_13065_),
    .B(_13064_),
    .X(_13202_));
 sky130_fd_sc_hd__nand2_1 _19922_ (.A(_11043_),
    .B(_11895_),
    .Y(_13203_));
 sky130_fd_sc_hd__and4_1 _19923_ (.A(_11174_),
    .B(_11903_),
    .C(_11889_),
    .D(_12020_),
    .X(_13204_));
 sky130_fd_sc_hd__a22o_1 _19924_ (.A1(_11903_),
    .A2(_11889_),
    .B1(_12020_),
    .B2(_11174_),
    .X(_13205_));
 sky130_fd_sc_hd__and2b_1 _19925_ (.A_N(_13204_),
    .B(_13205_),
    .X(_13206_));
 sky130_fd_sc_hd__xnor2_1 _19926_ (.A(_13203_),
    .B(_13206_),
    .Y(_13207_));
 sky130_fd_sc_hd__nand2_1 _19927_ (.A(_10852_),
    .B(\genblk1.pcpi_mul.rs2[21] ),
    .Y(_13208_));
 sky130_fd_sc_hd__and4_1 _19928_ (.A(_10848_),
    .B(_10745_),
    .C(_12327_),
    .D(_12464_),
    .X(_13209_));
 sky130_fd_sc_hd__a22oi_2 _19929_ (.A1(_10792_),
    .A2(_12322_),
    .B1(_12600_),
    .B2(_10696_),
    .Y(_13210_));
 sky130_fd_sc_hd__or3_1 _19930_ (.A(_13208_),
    .B(_13209_),
    .C(_13210_),
    .X(_13211_));
 sky130_fd_sc_hd__o21ai_1 _19931_ (.A1(_13209_),
    .A2(_13210_),
    .B1(_13208_),
    .Y(_13212_));
 sky130_fd_sc_hd__a21bo_1 _19932_ (.A1(_13075_),
    .A2(_13077_),
    .B1_N(_13076_),
    .X(_13213_));
 sky130_fd_sc_hd__nand3_1 _19933_ (.A(_13211_),
    .B(_13212_),
    .C(_13213_),
    .Y(_13214_));
 sky130_fd_sc_hd__a21o_1 _19934_ (.A1(_13211_),
    .A2(_13212_),
    .B1(_13213_),
    .X(_13215_));
 sky130_fd_sc_hd__nand3_2 _19935_ (.A(_13207_),
    .B(_13214_),
    .C(_13215_),
    .Y(_13216_));
 sky130_fd_sc_hd__a21o_1 _19936_ (.A1(_13214_),
    .A2(_13215_),
    .B1(_13207_),
    .X(_13217_));
 sky130_fd_sc_hd__nand3_4 _19937_ (.A(_13202_),
    .B(_13216_),
    .C(_13217_),
    .Y(_13218_));
 sky130_fd_sc_hd__a21o_1 _19938_ (.A1(_13216_),
    .A2(_13217_),
    .B1(_13202_),
    .X(_13219_));
 sky130_fd_sc_hd__nand3_2 _19939_ (.A(_13201_),
    .B(_13218_),
    .C(_13219_),
    .Y(_13220_));
 sky130_fd_sc_hd__a21o_1 _19940_ (.A1(_13218_),
    .A2(_13219_),
    .B1(_13201_),
    .X(_13221_));
 sky130_fd_sc_hd__or2b_1 _19941_ (.A(_13057_),
    .B_N(_13066_),
    .X(_13222_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19942_ (.A(\genblk1.pcpi_mul.rs2[28] ),
    .X(_13223_));
 sky130_fd_sc_hd__clkbuf_4 _19943_ (.A(_13223_),
    .X(_13224_));
 sky130_fd_sc_hd__a22o_1 _19944_ (.A1(_10636_),
    .A2(_13055_),
    .B1(_13224_),
    .B2(_10589_),
    .X(_13225_));
 sky130_fd_sc_hd__buf_2 _19945_ (.A(_13054_),
    .X(_13226_));
 sky130_fd_sc_hd__clkbuf_2 _19946_ (.A(\genblk1.pcpi_mul.rs2[28] ),
    .X(_13227_));
 sky130_fd_sc_hd__clkbuf_4 _19947_ (.A(_13227_),
    .X(_13228_));
 sky130_fd_sc_hd__clkbuf_4 _19948_ (.A(_13228_),
    .X(_13229_));
 sky130_fd_sc_hd__nand4_4 _19949_ (.A(_10589_),
    .B(_10596_),
    .C(_13226_),
    .D(_13229_),
    .Y(_13230_));
 sky130_fd_sc_hd__nand2_1 _19950_ (.A(_13225_),
    .B(_13230_),
    .Y(_13231_));
 sky130_fd_sc_hd__o21ba_1 _19951_ (.A1(_13058_),
    .A2(_13062_),
    .B1_N(_13059_),
    .X(_13232_));
 sky130_fd_sc_hd__nand2_1 _19952_ (.A(_10721_),
    .B(_12775_),
    .Y(_13233_));
 sky130_fd_sc_hd__and4_1 _19953_ (.A(_10752_),
    .B(_10648_),
    .C(_12909_),
    .D(\genblk1.pcpi_mul.rs2[26] ),
    .X(_13234_));
 sky130_fd_sc_hd__a22oi_2 _19954_ (.A1(_10717_),
    .A2(_12770_),
    .B1(_13061_),
    .B2(_10754_),
    .Y(_13235_));
 sky130_fd_sc_hd__nor2_1 _19955_ (.A(_13234_),
    .B(_13235_),
    .Y(_13236_));
 sky130_fd_sc_hd__xnor2_1 _19956_ (.A(_13233_),
    .B(_13236_),
    .Y(_13237_));
 sky130_fd_sc_hd__xnor2_1 _19957_ (.A(_13232_),
    .B(_13237_),
    .Y(_13238_));
 sky130_fd_sc_hd__xor2_2 _19958_ (.A(_13231_),
    .B(_13238_),
    .X(_13239_));
 sky130_fd_sc_hd__xor2_1 _19959_ (.A(_13222_),
    .B(_13239_),
    .X(_13240_));
 sky130_fd_sc_hd__nand3_1 _19960_ (.A(_13220_),
    .B(_13221_),
    .C(_13240_),
    .Y(_13241_));
 sky130_fd_sc_hd__a21o_1 _19961_ (.A1(_13220_),
    .A2(_13221_),
    .B1(_13240_),
    .X(_13242_));
 sky130_fd_sc_hd__nand3_1 _19962_ (.A(_13089_),
    .B(_13241_),
    .C(_13242_),
    .Y(_13243_));
 sky130_fd_sc_hd__a21o_1 _19963_ (.A1(_13241_),
    .A2(_13242_),
    .B1(_13089_),
    .X(_13244_));
 sky130_fd_sc_hd__and4_2 _19964_ (.A(_13199_),
    .B(_13200_),
    .C(_13243_),
    .D(_13244_),
    .X(_13245_));
 sky130_fd_sc_hd__a22oi_2 _19965_ (.A1(_13199_),
    .A2(_13200_),
    .B1(_13243_),
    .B2(_13244_),
    .Y(_13246_));
 sky130_fd_sc_hd__a211o_1 _19966_ (.A1(_13091_),
    .A2(_13093_),
    .B1(_13245_),
    .C1(_13246_),
    .X(_13247_));
 sky130_fd_sc_hd__o211ai_2 _19967_ (.A1(_13245_),
    .A2(_13246_),
    .B1(_13091_),
    .C1(_13093_),
    .Y(_13248_));
 sky130_fd_sc_hd__nand4_1 _19968_ (.A(_13163_),
    .B(_13164_),
    .C(_13247_),
    .D(_13248_),
    .Y(_13249_));
 sky130_fd_sc_hd__a22o_1 _19969_ (.A1(_13163_),
    .A2(_13164_),
    .B1(_13247_),
    .B2(_13248_),
    .X(_13250_));
 sky130_fd_sc_hd__o211a_1 _19970_ (.A1(_13095_),
    .A2(net417),
    .B1(_13249_),
    .C1(_13250_),
    .X(_13251_));
 sky130_fd_sc_hd__a211oi_1 _19971_ (.A1(_13249_),
    .A2(_13250_),
    .B1(_13095_),
    .C1(net417),
    .Y(_13252_));
 sky130_fd_sc_hd__or3_1 _19972_ (.A(_13116_),
    .B(_13251_),
    .C(_13252_),
    .X(_13253_));
 sky130_fd_sc_hd__o21ai_1 _19973_ (.A1(_13251_),
    .A2(_13252_),
    .B1(_13116_),
    .Y(_13254_));
 sky130_fd_sc_hd__o211a_1 _19974_ (.A1(_13099_),
    .A2(_13113_),
    .B1(_13253_),
    .C1(_13254_),
    .X(_13255_));
 sky130_fd_sc_hd__a211oi_1 _19975_ (.A1(_13253_),
    .A2(_13254_),
    .B1(_13099_),
    .C1(_13113_),
    .Y(_13256_));
 sky130_fd_sc_hd__nor3_1 _19976_ (.A(_13112_),
    .B(_13255_),
    .C(_13256_),
    .Y(_13257_));
 sky130_fd_sc_hd__o21a_1 _19977_ (.A1(_13255_),
    .A2(_13256_),
    .B1(_13112_),
    .X(_13258_));
 sky130_fd_sc_hd__or2_2 _19978_ (.A(_13257_),
    .B(_13258_),
    .X(_13259_));
 sky130_fd_sc_hd__and2b_1 _19979_ (.A_N(_13103_),
    .B(_13105_),
    .X(_13260_));
 sky130_fd_sc_hd__xnor2_2 _19980_ (.A(_13259_),
    .B(_13260_),
    .Y(_13261_));
 sky130_fd_sc_hd__or4_1 _19981_ (.A(_12953_),
    .B(_12954_),
    .C(_13108_),
    .D(_13109_),
    .X(_13262_));
 sky130_fd_sc_hd__a211o_1 _19982_ (.A1(_13105_),
    .A2(_13106_),
    .B1(_12949_),
    .C1(_13107_),
    .X(_13263_));
 sky130_fd_sc_hd__a21oi_1 _19983_ (.A1(_12953_),
    .A2(_13263_),
    .B1(_13109_),
    .Y(_13264_));
 sky130_fd_sc_hd__o21a_1 _19984_ (.A1(_12958_),
    .A2(_13262_),
    .B1(_13264_),
    .X(_13265_));
 sky130_fd_sc_hd__xor2_1 _19985_ (.A(_13261_),
    .B(_13265_),
    .X(_00074_));
 sky130_fd_sc_hd__o21ai_1 _19986_ (.A1(_12990_),
    .A2(_12992_),
    .B1(_13114_),
    .Y(_13266_));
 sky130_fd_sc_hd__nor3_1 _19987_ (.A(_13116_),
    .B(_13251_),
    .C(_13252_),
    .Y(_13267_));
 sky130_fd_sc_hd__nor2_1 _19988_ (.A(_13137_),
    .B(_13139_),
    .Y(_13268_));
 sky130_fd_sc_hd__a21o_1 _19989_ (.A1(_13161_),
    .A2(_13163_),
    .B1(_13268_),
    .X(_13269_));
 sky130_fd_sc_hd__nand3_1 _19990_ (.A(_13161_),
    .B(_13163_),
    .C(_13268_),
    .Y(_13270_));
 sky130_fd_sc_hd__nand2_1 _19991_ (.A(_13269_),
    .B(_13270_),
    .Y(_13271_));
 sky130_vsdinv _19992_ (.A(_13247_),
    .Y(_13272_));
 sky130_fd_sc_hd__and4_1 _19993_ (.A(_13163_),
    .B(_13164_),
    .C(_13247_),
    .D(_13248_),
    .X(_13273_));
 sky130_fd_sc_hd__nand2_1 _19994_ (.A(_13157_),
    .B(_13159_),
    .Y(_13274_));
 sky130_fd_sc_hd__a211o_1 _19995_ (.A1(_13085_),
    .A2(_13087_),
    .B1(net366),
    .C1(_13196_),
    .X(_13275_));
 sky130_fd_sc_hd__or2_1 _19996_ (.A(_12972_),
    .B(_13122_),
    .X(_13276_));
 sky130_fd_sc_hd__a211o_1 _19997_ (.A1(_12974_),
    .A2(_13121_),
    .B1(_13126_),
    .C1(_13123_),
    .X(_13277_));
 sky130_fd_sc_hd__or2b_1 _19998_ (.A(_13134_),
    .B_N(_13133_),
    .X(_13278_));
 sky130_fd_sc_hd__nand2_1 _19999_ (.A(_13127_),
    .B(_13135_),
    .Y(_13279_));
 sky130_fd_sc_hd__nand2_1 _20000_ (.A(_10747_),
    .B(_13128_),
    .Y(_13280_));
 sky130_fd_sc_hd__clkbuf_4 _20001_ (.A(\genblk1.pcpi_mul.rs1[28] ),
    .X(_13281_));
 sky130_fd_sc_hd__nand2_2 _20002_ (.A(_10611_),
    .B(_13281_),
    .Y(_13282_));
 sky130_fd_sc_hd__nor2_1 _20003_ (.A(_13121_),
    .B(_13282_),
    .Y(_13283_));
 sky130_fd_sc_hd__a21oi_1 _20004_ (.A1(_13122_),
    .A2(_13280_),
    .B1(_13283_),
    .Y(_13284_));
 sky130_fd_sc_hd__clkbuf_2 _20005_ (.A(_12973_),
    .X(_13285_));
 sky130_fd_sc_hd__buf_4 _20006_ (.A(_13285_),
    .X(_13286_));
 sky130_fd_sc_hd__nand2_2 _20007_ (.A(_11704_),
    .B(_13286_),
    .Y(_13287_));
 sky130_fd_sc_hd__xnor2_1 _20008_ (.A(_13284_),
    .B(_13287_),
    .Y(_13288_));
 sky130_fd_sc_hd__and4_1 _20009_ (.A(_10700_),
    .B(_10803_),
    .C(_12688_),
    .D(\genblk1.pcpi_mul.rs1[25] ),
    .X(_13289_));
 sky130_fd_sc_hd__a22oi_2 _20010_ (.A1(_11711_),
    .A2(_12688_),
    .B1(_12700_),
    .B2(_10671_),
    .Y(_13290_));
 sky130_fd_sc_hd__nor2_1 _20011_ (.A(_13289_),
    .B(_13290_),
    .Y(_13291_));
 sky130_fd_sc_hd__clkbuf_4 _20012_ (.A(\genblk1.pcpi_mul.rs1[29] ),
    .X(_13292_));
 sky130_fd_sc_hd__nand2_1 _20013_ (.A(_10583_),
    .B(_13292_),
    .Y(_13293_));
 sky130_fd_sc_hd__xnor2_1 _20014_ (.A(_13291_),
    .B(_13293_),
    .Y(_13294_));
 sky130_fd_sc_hd__o21ba_1 _20015_ (.A1(_13129_),
    .A2(_13131_),
    .B1_N(_13130_),
    .X(_13295_));
 sky130_fd_sc_hd__xnor2_1 _20016_ (.A(_13294_),
    .B(_13295_),
    .Y(_13296_));
 sky130_fd_sc_hd__xnor2_1 _20017_ (.A(_13288_),
    .B(_13296_),
    .Y(_13297_));
 sky130_fd_sc_hd__a21oi_1 _20018_ (.A1(_13278_),
    .A2(_13279_),
    .B1(_13297_),
    .Y(_13298_));
 sky130_fd_sc_hd__and3_1 _20019_ (.A(_13278_),
    .B(_13279_),
    .C(_13297_),
    .X(_13299_));
 sky130_fd_sc_hd__a211oi_2 _20020_ (.A1(_13276_),
    .A2(_13277_),
    .B1(_13298_),
    .C1(_13299_),
    .Y(_13300_));
 sky130_fd_sc_hd__o211a_1 _20021_ (.A1(_13298_),
    .A2(_13299_),
    .B1(_13276_),
    .C1(_13277_),
    .X(_13301_));
 sky130_fd_sc_hd__nand3_1 _20022_ (.A(_13141_),
    .B(_13151_),
    .C(_13152_),
    .Y(_13302_));
 sky130_fd_sc_hd__a21o_1 _20023_ (.A1(_13170_),
    .A2(_13178_),
    .B1(_13177_),
    .X(_13303_));
 sky130_fd_sc_hd__nand2_1 _20024_ (.A(_13145_),
    .B(_13147_),
    .Y(_13304_));
 sky130_fd_sc_hd__clkbuf_4 _20025_ (.A(_12069_),
    .X(_13305_));
 sky130_fd_sc_hd__a31o_1 _20026_ (.A1(_10960_),
    .A2(_13305_),
    .A3(_13168_),
    .B1(_13167_),
    .X(_13306_));
 sky130_fd_sc_hd__a22o_1 _20027_ (.A1(_11195_),
    .A2(_12273_),
    .B1(_12281_),
    .B2(_12172_),
    .X(_13307_));
 sky130_fd_sc_hd__nand4_2 _20028_ (.A(_10997_),
    .B(_11085_),
    .C(_12273_),
    .D(_12281_),
    .Y(_13308_));
 sky130_fd_sc_hd__a22o_1 _20029_ (.A1(_10993_),
    .A2(_12538_),
    .B1(_13307_),
    .B2(_13308_),
    .X(_13309_));
 sky130_fd_sc_hd__nand4_2 _20030_ (.A(_11508_),
    .B(_12416_),
    .C(_13307_),
    .D(_13308_),
    .Y(_13310_));
 sky130_fd_sc_hd__nand3_2 _20031_ (.A(_13306_),
    .B(_13309_),
    .C(_13310_),
    .Y(_13311_));
 sky130_fd_sc_hd__a21o_1 _20032_ (.A1(_13309_),
    .A2(_13310_),
    .B1(_13306_),
    .X(_13312_));
 sky130_fd_sc_hd__nand3_1 _20033_ (.A(_13304_),
    .B(_13311_),
    .C(_13312_),
    .Y(_13313_));
 sky130_fd_sc_hd__a21o_1 _20034_ (.A1(_13311_),
    .A2(_13312_),
    .B1(_13304_),
    .X(_13314_));
 sky130_fd_sc_hd__and3_1 _20035_ (.A(_13303_),
    .B(_13313_),
    .C(_13314_),
    .X(_13315_));
 sky130_fd_sc_hd__a21oi_1 _20036_ (.A1(_13313_),
    .A2(_13314_),
    .B1(_13303_),
    .Y(_13316_));
 sky130_fd_sc_hd__a211oi_2 _20037_ (.A1(_13149_),
    .A2(_13151_),
    .B1(_13315_),
    .C1(_13316_),
    .Y(_13317_));
 sky130_fd_sc_hd__o211a_1 _20038_ (.A1(_13315_),
    .A2(_13316_),
    .B1(_13149_),
    .C1(_13151_),
    .X(_13318_));
 sky130_fd_sc_hd__a211oi_2 _20039_ (.A1(_13302_),
    .A2(_13155_),
    .B1(_13317_),
    .C1(_13318_),
    .Y(_13319_));
 sky130_fd_sc_hd__o211a_1 _20040_ (.A1(_13317_),
    .A2(_13318_),
    .B1(_13302_),
    .C1(_13155_),
    .X(_13320_));
 sky130_fd_sc_hd__nor4_2 _20041_ (.A(_13300_),
    .B(_13301_),
    .C(_13319_),
    .D(_13320_),
    .Y(_13321_));
 sky130_fd_sc_hd__o22a_1 _20042_ (.A1(_13300_),
    .A2(_13301_),
    .B1(_13319_),
    .B2(_13320_),
    .X(_13322_));
 sky130_fd_sc_hd__a211o_1 _20043_ (.A1(_13275_),
    .A2(_13199_),
    .B1(net362),
    .C1(_13322_),
    .X(_13323_));
 sky130_fd_sc_hd__o211ai_2 _20044_ (.A1(net362),
    .A2(_13322_),
    .B1(_13275_),
    .C1(_13199_),
    .Y(_13324_));
 sky130_fd_sc_hd__nand3_2 _20045_ (.A(_13274_),
    .B(_13323_),
    .C(_13324_),
    .Y(_13325_));
 sky130_fd_sc_hd__a21o_1 _20046_ (.A1(_13323_),
    .A2(_13324_),
    .B1(_13274_),
    .X(_13326_));
 sky130_fd_sc_hd__and3_1 _20047_ (.A(_13089_),
    .B(_13241_),
    .C(_13242_),
    .X(_13327_));
 sky130_vsdinv _20048_ (.A(_13193_),
    .Y(_13328_));
 sky130_vsdinv _20049_ (.A(_13195_),
    .Y(_13329_));
 sky130_fd_sc_hd__nand2_1 _20050_ (.A(_10892_),
    .B(_12079_),
    .Y(_13330_));
 sky130_fd_sc_hd__and4_1 _20051_ (.A(_10955_),
    .B(_11106_),
    .C(_11945_),
    .D(_11957_),
    .X(_13331_));
 sky130_fd_sc_hd__a22o_1 _20052_ (.A1(_11110_),
    .A2(_11945_),
    .B1(_11957_),
    .B2(_10955_),
    .X(_13332_));
 sky130_fd_sc_hd__and2b_1 _20053_ (.A_N(_13331_),
    .B(_13332_),
    .X(_13333_));
 sky130_fd_sc_hd__xnor2_1 _20054_ (.A(_13330_),
    .B(_13333_),
    .Y(_13334_));
 sky130_fd_sc_hd__nand2_1 _20055_ (.A(_11349_),
    .B(_11818_),
    .Y(_13335_));
 sky130_fd_sc_hd__and4_1 _20056_ (.A(_11240_),
    .B(_11457_),
    .C(_11588_),
    .D(_11697_),
    .X(_13336_));
 sky130_fd_sc_hd__a22oi_2 _20057_ (.A1(_11353_),
    .A2(_11488_),
    .B1(_11597_),
    .B2(_11795_),
    .Y(_13337_));
 sky130_fd_sc_hd__or3_1 _20058_ (.A(_13335_),
    .B(_13336_),
    .C(_13337_),
    .X(_13338_));
 sky130_fd_sc_hd__o21ai_1 _20059_ (.A1(_13336_),
    .A2(_13337_),
    .B1(_13335_),
    .Y(_13339_));
 sky130_fd_sc_hd__o21bai_1 _20060_ (.A1(_13171_),
    .A2(_13173_),
    .B1_N(_13172_),
    .Y(_13340_));
 sky130_fd_sc_hd__and3_1 _20061_ (.A(_13338_),
    .B(_13339_),
    .C(_13340_),
    .X(_13341_));
 sky130_fd_sc_hd__a21o_1 _20062_ (.A1(_13338_),
    .A2(_13339_),
    .B1(_13340_),
    .X(_13342_));
 sky130_fd_sc_hd__and2b_1 _20063_ (.A_N(_13341_),
    .B(_13342_),
    .X(_13343_));
 sky130_fd_sc_hd__xnor2_1 _20064_ (.A(_13334_),
    .B(_13343_),
    .Y(_13344_));
 sky130_fd_sc_hd__nand2_1 _20065_ (.A(_13184_),
    .B(_13186_),
    .Y(_13345_));
 sky130_fd_sc_hd__a31o_1 _20066_ (.A1(_11269_),
    .A2(_11894_),
    .A3(_13205_),
    .B1(_13204_),
    .X(_13346_));
 sky130_fd_sc_hd__nand4_2 _20067_ (.A(_11260_),
    .B(_11276_),
    .C(_11662_),
    .D(_11924_),
    .Y(_13347_));
 sky130_fd_sc_hd__a22o_1 _20068_ (.A1(_11371_),
    .A2(_11922_),
    .B1(_11780_),
    .B2(_12098_),
    .X(_13348_));
 sky130_fd_sc_hd__nand4_2 _20069_ (.A(_12561_),
    .B(_11559_),
    .C(_13347_),
    .D(_13348_),
    .Y(_13349_));
 sky130_fd_sc_hd__a22o_1 _20070_ (.A1(_11834_),
    .A2(_11443_),
    .B1(_13347_),
    .B2(_13348_),
    .X(_13350_));
 sky130_fd_sc_hd__nand3_1 _20071_ (.A(_13346_),
    .B(_13349_),
    .C(_13350_),
    .Y(_13351_));
 sky130_fd_sc_hd__a21o_1 _20072_ (.A1(_13349_),
    .A2(_13350_),
    .B1(_13346_),
    .X(_13352_));
 sky130_fd_sc_hd__nand3_1 _20073_ (.A(_13345_),
    .B(_13351_),
    .C(_13352_),
    .Y(_13353_));
 sky130_fd_sc_hd__a21o_1 _20074_ (.A1(_13351_),
    .A2(_13352_),
    .B1(_13345_),
    .X(_13354_));
 sky130_fd_sc_hd__a21bo_1 _20075_ (.A1(_13181_),
    .A2(_13189_),
    .B1_N(_13188_),
    .X(_13355_));
 sky130_fd_sc_hd__and3_1 _20076_ (.A(_13353_),
    .B(_13354_),
    .C(_13355_),
    .X(_13356_));
 sky130_fd_sc_hd__a21oi_1 _20077_ (.A1(_13353_),
    .A2(_13354_),
    .B1(_13355_),
    .Y(_13357_));
 sky130_fd_sc_hd__nor3_2 _20078_ (.A(_13344_),
    .B(_13356_),
    .C(_13357_),
    .Y(_13358_));
 sky130_fd_sc_hd__o21a_1 _20079_ (.A1(_13356_),
    .A2(_13357_),
    .B1(_13344_),
    .X(_13359_));
 sky130_fd_sc_hd__a211oi_4 _20080_ (.A1(_13218_),
    .A2(_13220_),
    .B1(_13358_),
    .C1(_13359_),
    .Y(_13360_));
 sky130_fd_sc_hd__o211a_1 _20081_ (.A1(_13358_),
    .A2(_13359_),
    .B1(_13218_),
    .C1(_13220_),
    .X(_13361_));
 sky130_fd_sc_hd__a211oi_2 _20082_ (.A1(_13328_),
    .A2(_13329_),
    .B1(_13360_),
    .C1(_13361_),
    .Y(_13362_));
 sky130_fd_sc_hd__o211a_1 _20083_ (.A1(_13360_),
    .A2(_13361_),
    .B1(_13328_),
    .C1(_13329_),
    .X(_13363_));
 sky130_fd_sc_hd__nor2_1 _20084_ (.A(_13222_),
    .B(_13239_),
    .Y(_13364_));
 sky130_fd_sc_hd__and3_1 _20085_ (.A(_13220_),
    .B(_13221_),
    .C(_13240_),
    .X(_13365_));
 sky130_fd_sc_hd__nand2_1 _20086_ (.A(_13214_),
    .B(_13216_),
    .Y(_13366_));
 sky130_fd_sc_hd__and2b_1 _20087_ (.A_N(_13232_),
    .B(_13237_),
    .X(_13367_));
 sky130_fd_sc_hd__nand2_1 _20088_ (.A(_11056_),
    .B(_11895_),
    .Y(_13368_));
 sky130_fd_sc_hd__and4_1 _20089_ (.A(_10919_),
    .B(_11268_),
    .C(_11889_),
    .D(_12233_),
    .X(_13369_));
 sky130_fd_sc_hd__a22o_1 _20090_ (.A1(_11268_),
    .A2(_12235_),
    .B1(_12233_),
    .B2(_10919_),
    .X(_13370_));
 sky130_fd_sc_hd__and2b_1 _20091_ (.A_N(_13369_),
    .B(_13370_),
    .X(_13371_));
 sky130_fd_sc_hd__xnor2_1 _20092_ (.A(_13368_),
    .B(_13371_),
    .Y(_13372_));
 sky130_fd_sc_hd__and2_1 _20093_ (.A(_10967_),
    .B(\genblk1.pcpi_mul.rs2[21] ),
    .X(_13373_));
 sky130_fd_sc_hd__clkbuf_2 _20094_ (.A(_12600_),
    .X(_13374_));
 sky130_fd_sc_hd__nand4_4 _20095_ (.A(_10757_),
    .B(_11062_),
    .C(_12328_),
    .D(_13374_),
    .Y(_13375_));
 sky130_fd_sc_hd__buf_2 _20096_ (.A(_12464_),
    .X(_13376_));
 sky130_fd_sc_hd__a22o_1 _20097_ (.A1(_10805_),
    .A2(_12322_),
    .B1(_13376_),
    .B2(_11301_),
    .X(_13377_));
 sky130_fd_sc_hd__nand3_1 _20098_ (.A(_13373_),
    .B(_13375_),
    .C(_13377_),
    .Y(_13378_));
 sky130_fd_sc_hd__a21o_1 _20099_ (.A1(_13375_),
    .A2(_13377_),
    .B1(_13373_),
    .X(_13379_));
 sky130_fd_sc_hd__o21bai_1 _20100_ (.A1(_13208_),
    .A2(_13210_),
    .B1_N(_13209_),
    .Y(_13380_));
 sky130_fd_sc_hd__nand3_2 _20101_ (.A(_13378_),
    .B(_13379_),
    .C(_13380_),
    .Y(_13381_));
 sky130_fd_sc_hd__a21o_1 _20102_ (.A1(_13378_),
    .A2(_13379_),
    .B1(_13380_),
    .X(_13382_));
 sky130_fd_sc_hd__nand3_2 _20103_ (.A(_13372_),
    .B(_13381_),
    .C(_13382_),
    .Y(_13383_));
 sky130_fd_sc_hd__a21o_1 _20104_ (.A1(_13381_),
    .A2(_13382_),
    .B1(_13372_),
    .X(_13384_));
 sky130_fd_sc_hd__nand3_4 _20105_ (.A(_13367_),
    .B(_13383_),
    .C(_13384_),
    .Y(_13385_));
 sky130_fd_sc_hd__a21o_1 _20106_ (.A1(_13383_),
    .A2(_13384_),
    .B1(_13367_),
    .X(_13386_));
 sky130_fd_sc_hd__nand3_4 _20107_ (.A(_13366_),
    .B(_13385_),
    .C(_13386_),
    .Y(_13387_));
 sky130_fd_sc_hd__a21o_1 _20108_ (.A1(_13385_),
    .A2(_13386_),
    .B1(_13366_),
    .X(_13388_));
 sky130_fd_sc_hd__nand2_1 _20109_ (.A(_10630_),
    .B(_13055_),
    .Y(_13389_));
 sky130_fd_sc_hd__and4_1 _20110_ (.A(_10587_),
    .B(_10786_),
    .C(_13227_),
    .D(\genblk1.pcpi_mul.rs2[29] ),
    .X(_13390_));
 sky130_fd_sc_hd__a22o_1 _20111_ (.A1(_10705_),
    .A2(_13227_),
    .B1(\genblk1.pcpi_mul.rs2[29] ),
    .B2(_10587_),
    .X(_13391_));
 sky130_fd_sc_hd__and2b_1 _20112_ (.A_N(_13390_),
    .B(_13391_),
    .X(_13392_));
 sky130_fd_sc_hd__xnor2_1 _20113_ (.A(_13389_),
    .B(_13392_),
    .Y(_13393_));
 sky130_fd_sc_hd__a31o_1 _20114_ (.A1(_10666_),
    .A2(_12584_),
    .A3(_13236_),
    .B1(_13234_),
    .X(_13394_));
 sky130_fd_sc_hd__and4_1 _20115_ (.A(_10710_),
    .B(_10705_),
    .C(\genblk1.pcpi_mul.rs2[27] ),
    .D(_13227_),
    .X(_13395_));
 sky130_fd_sc_hd__nand4_2 _20116_ (.A(_10648_),
    .B(_10741_),
    .C(_12909_),
    .D(_12910_),
    .Y(_13396_));
 sky130_fd_sc_hd__a22o_1 _20117_ (.A1(_10664_),
    .A2(_12909_),
    .B1(\genblk1.pcpi_mul.rs2[26] ),
    .B2(_10800_),
    .X(_13397_));
 sky130_fd_sc_hd__nand4_1 _20118_ (.A(_10697_),
    .B(_12775_),
    .C(_13396_),
    .D(_13397_),
    .Y(_13398_));
 sky130_fd_sc_hd__a22o_1 _20119_ (.A1(_10746_),
    .A2(\genblk1.pcpi_mul.rs2[24] ),
    .B1(_13396_),
    .B2(_13397_),
    .X(_13399_));
 sky130_fd_sc_hd__nand3_1 _20120_ (.A(_13395_),
    .B(_13398_),
    .C(_13399_),
    .Y(_13400_));
 sky130_fd_sc_hd__a21o_1 _20121_ (.A1(_13398_),
    .A2(_13399_),
    .B1(_13395_),
    .X(_13401_));
 sky130_fd_sc_hd__nand3_1 _20122_ (.A(_13394_),
    .B(_13400_),
    .C(_13401_),
    .Y(_13402_));
 sky130_fd_sc_hd__a21o_1 _20123_ (.A1(_13400_),
    .A2(_13401_),
    .B1(_13394_),
    .X(_13403_));
 sky130_fd_sc_hd__and3_1 _20124_ (.A(_13393_),
    .B(_13402_),
    .C(_13403_),
    .X(_13404_));
 sky130_fd_sc_hd__a21oi_1 _20125_ (.A1(_13402_),
    .A2(_13403_),
    .B1(_13393_),
    .Y(_13405_));
 sky130_fd_sc_hd__and3_1 _20126_ (.A(_13225_),
    .B(_13230_),
    .C(_13238_),
    .X(_13406_));
 sky130_fd_sc_hd__or3b_4 _20127_ (.A(_13404_),
    .B(_13405_),
    .C_N(_13406_),
    .X(_13407_));
 sky130_fd_sc_hd__o21bai_2 _20128_ (.A1(_13404_),
    .A2(_13405_),
    .B1_N(_13406_),
    .Y(_13408_));
 sky130_fd_sc_hd__nand4_4 _20129_ (.A(_13387_),
    .B(_13388_),
    .C(_13407_),
    .D(_13408_),
    .Y(_13409_));
 sky130_fd_sc_hd__a22o_1 _20130_ (.A1(_13387_),
    .A2(_13388_),
    .B1(_13407_),
    .B2(_13408_),
    .X(_13410_));
 sky130_fd_sc_hd__o211ai_2 _20131_ (.A1(_13364_),
    .A2(_13365_),
    .B1(_13409_),
    .C1(_13410_),
    .Y(_13411_));
 sky130_fd_sc_hd__a211o_1 _20132_ (.A1(_13409_),
    .A2(_13410_),
    .B1(_13364_),
    .C1(_13365_),
    .X(_13412_));
 sky130_fd_sc_hd__or4bb_4 _20133_ (.A(_13362_),
    .B(_13363_),
    .C_N(_13411_),
    .D_N(_13412_),
    .X(_13413_));
 sky130_fd_sc_hd__a2bb2o_1 _20134_ (.A1_N(_13362_),
    .A2_N(_13363_),
    .B1(_13411_),
    .B2(_13412_),
    .X(_13414_));
 sky130_fd_sc_hd__o211ai_4 _20135_ (.A1(_13327_),
    .A2(_13245_),
    .B1(_13413_),
    .C1(_13414_),
    .Y(_13415_));
 sky130_fd_sc_hd__a211o_1 _20136_ (.A1(_13413_),
    .A2(_13414_),
    .B1(_13327_),
    .C1(_13245_),
    .X(_13416_));
 sky130_fd_sc_hd__nand4_2 _20137_ (.A(_13325_),
    .B(_13326_),
    .C(_13415_),
    .D(_13416_),
    .Y(_13417_));
 sky130_fd_sc_hd__a22o_1 _20138_ (.A1(_13325_),
    .A2(_13326_),
    .B1(_13415_),
    .B2(_13416_),
    .X(_13418_));
 sky130_fd_sc_hd__o211a_1 _20139_ (.A1(_13272_),
    .A2(_13273_),
    .B1(_13417_),
    .C1(_13418_),
    .X(_13419_));
 sky130_fd_sc_hd__a211oi_1 _20140_ (.A1(_13417_),
    .A2(_13418_),
    .B1(_13272_),
    .C1(_13273_),
    .Y(_13420_));
 sky130_fd_sc_hd__or3_1 _20141_ (.A(_13271_),
    .B(_13419_),
    .C(_13420_),
    .X(_13421_));
 sky130_fd_sc_hd__o21ai_1 _20142_ (.A1(_13419_),
    .A2(_13420_),
    .B1(_13271_),
    .Y(_13422_));
 sky130_fd_sc_hd__o211a_1 _20143_ (.A1(_13251_),
    .A2(_13267_),
    .B1(_13421_),
    .C1(_13422_),
    .X(_13423_));
 sky130_fd_sc_hd__a211oi_1 _20144_ (.A1(_13421_),
    .A2(_13422_),
    .B1(_13251_),
    .C1(_13267_),
    .Y(_13424_));
 sky130_fd_sc_hd__or3_1 _20145_ (.A(_13266_),
    .B(_13423_),
    .C(_13424_),
    .X(_13425_));
 sky130_fd_sc_hd__o21ai_1 _20146_ (.A1(_13423_),
    .A2(_13424_),
    .B1(_13266_),
    .Y(_13426_));
 sky130_fd_sc_hd__o211a_1 _20147_ (.A1(_13255_),
    .A2(_13257_),
    .B1(_13425_),
    .C1(_13426_),
    .X(_13427_));
 sky130_fd_sc_hd__a211oi_2 _20148_ (.A1(_13425_),
    .A2(_13426_),
    .B1(_13255_),
    .C1(_13257_),
    .Y(_13428_));
 sky130_fd_sc_hd__or2_1 _20149_ (.A(_13427_),
    .B(_13428_),
    .X(_13429_));
 sky130_fd_sc_hd__or2_1 _20150_ (.A(_13259_),
    .B(_13260_),
    .X(_13430_));
 sky130_fd_sc_hd__o21ai_1 _20151_ (.A1(_13261_),
    .A2(_13265_),
    .B1(_13430_),
    .Y(_13431_));
 sky130_fd_sc_hd__xnor2_1 _20152_ (.A(_13429_),
    .B(_13431_),
    .Y(_00075_));
 sky130_fd_sc_hd__nor3_1 _20153_ (.A(_13271_),
    .B(_13419_),
    .C(_13420_),
    .Y(_13432_));
 sky130_fd_sc_hd__nor2_1 _20154_ (.A(_13298_),
    .B(_13300_),
    .Y(_13433_));
 sky130_fd_sc_hd__a21o_1 _20155_ (.A1(_13323_),
    .A2(_13325_),
    .B1(_13433_),
    .X(_13434_));
 sky130_fd_sc_hd__nand3_1 _20156_ (.A(_13323_),
    .B(_13325_),
    .C(_13433_),
    .Y(_13435_));
 sky130_fd_sc_hd__nand2_1 _20157_ (.A(_13434_),
    .B(_13435_),
    .Y(_13436_));
 sky130_fd_sc_hd__or2_1 _20158_ (.A(_13121_),
    .B(_13282_),
    .X(_13437_));
 sky130_fd_sc_hd__a211o_1 _20159_ (.A1(_13122_),
    .A2(_13280_),
    .B1(_13287_),
    .C1(_13283_),
    .X(_13438_));
 sky130_fd_sc_hd__or2b_1 _20160_ (.A(_13295_),
    .B_N(_13294_),
    .X(_13439_));
 sky130_fd_sc_hd__nand2_1 _20161_ (.A(_13288_),
    .B(_13296_),
    .Y(_13440_));
 sky130_fd_sc_hd__nand2_1 _20162_ (.A(_10600_),
    .B(_13292_),
    .Y(_13441_));
 sky130_fd_sc_hd__nand2_4 _20163_ (.A(_10740_),
    .B(\genblk1.pcpi_mul.rs1[29] ),
    .Y(_13442_));
 sky130_fd_sc_hd__nor2_1 _20164_ (.A(_13280_),
    .B(_13442_),
    .Y(_13443_));
 sky130_fd_sc_hd__a21oi_1 _20165_ (.A1(_13282_),
    .A2(_13441_),
    .B1(_13443_),
    .Y(_13444_));
 sky130_fd_sc_hd__clkbuf_2 _20166_ (.A(\genblk1.pcpi_mul.rs1[27] ),
    .X(_13445_));
 sky130_fd_sc_hd__clkbuf_4 _20167_ (.A(_13445_),
    .X(_13446_));
 sky130_fd_sc_hd__nand2_2 _20168_ (.A(_10644_),
    .B(_13446_),
    .Y(_13447_));
 sky130_fd_sc_hd__xnor2_1 _20169_ (.A(_13444_),
    .B(_13447_),
    .Y(_13448_));
 sky130_fd_sc_hd__a22oi_2 _20170_ (.A1(_10803_),
    .A2(\genblk1.pcpi_mul.rs1[25] ),
    .B1(\genblk1.pcpi_mul.rs1[26] ),
    .B2(_10700_),
    .Y(_13449_));
 sky130_fd_sc_hd__and4_1 _20171_ (.A(_10802_),
    .B(_10916_),
    .C(\genblk1.pcpi_mul.rs1[25] ),
    .D(\genblk1.pcpi_mul.rs1[26] ),
    .X(_13450_));
 sky130_fd_sc_hd__nor2_1 _20172_ (.A(_13449_),
    .B(_13450_),
    .Y(_13451_));
 sky130_fd_sc_hd__nand2_1 _20173_ (.A(_10583_),
    .B(\genblk1.pcpi_mul.rs1[30] ),
    .Y(_13452_));
 sky130_fd_sc_hd__xnor2_1 _20174_ (.A(_13451_),
    .B(_13452_),
    .Y(_13453_));
 sky130_fd_sc_hd__o21ba_1 _20175_ (.A1(_13290_),
    .A2(_13293_),
    .B1_N(_13289_),
    .X(_13454_));
 sky130_fd_sc_hd__xnor2_1 _20176_ (.A(_13453_),
    .B(_13454_),
    .Y(_13455_));
 sky130_fd_sc_hd__xnor2_1 _20177_ (.A(_13448_),
    .B(_13455_),
    .Y(_13456_));
 sky130_fd_sc_hd__a21oi_2 _20178_ (.A1(_13439_),
    .A2(_13440_),
    .B1(_13456_),
    .Y(_13457_));
 sky130_fd_sc_hd__and3_1 _20179_ (.A(_13439_),
    .B(_13440_),
    .C(_13456_),
    .X(_13458_));
 sky130_fd_sc_hd__a211oi_2 _20180_ (.A1(_13437_),
    .A2(_13438_),
    .B1(_13457_),
    .C1(_13458_),
    .Y(_13459_));
 sky130_fd_sc_hd__o211a_1 _20181_ (.A1(_13457_),
    .A2(_13458_),
    .B1(_13437_),
    .C1(_13438_),
    .X(_13460_));
 sky130_fd_sc_hd__a21o_1 _20182_ (.A1(_13334_),
    .A2(_13342_),
    .B1(_13341_),
    .X(_13461_));
 sky130_fd_sc_hd__nand2_1 _20183_ (.A(_13308_),
    .B(_13310_),
    .Y(_13462_));
 sky130_fd_sc_hd__a31o_1 _20184_ (.A1(_11189_),
    .A2(_12147_),
    .A3(_13332_),
    .B1(_13331_),
    .X(_13463_));
 sky130_fd_sc_hd__a22o_1 _20185_ (.A1(_11195_),
    .A2(\genblk1.pcpi_mul.rs1[22] ),
    .B1(\genblk1.pcpi_mul.rs1[23] ),
    .B2(_12172_),
    .X(_13464_));
 sky130_fd_sc_hd__nand4_2 _20186_ (.A(_10997_),
    .B(_11195_),
    .C(_12281_),
    .D(_12537_),
    .Y(_13465_));
 sky130_fd_sc_hd__a22o_1 _20187_ (.A1(_10993_),
    .A2(_12690_),
    .B1(_13464_),
    .B2(_13465_),
    .X(_13466_));
 sky130_fd_sc_hd__nand4_2 _20188_ (.A(_10736_),
    .B(_12690_),
    .C(_13464_),
    .D(_13465_),
    .Y(_13467_));
 sky130_fd_sc_hd__nand3_2 _20189_ (.A(_13463_),
    .B(_13466_),
    .C(_13467_),
    .Y(_13468_));
 sky130_fd_sc_hd__a21o_1 _20190_ (.A1(_13466_),
    .A2(_13467_),
    .B1(_13463_),
    .X(_13469_));
 sky130_fd_sc_hd__nand3_2 _20191_ (.A(_13462_),
    .B(_13468_),
    .C(_13469_),
    .Y(_13470_));
 sky130_fd_sc_hd__a21o_1 _20192_ (.A1(_13468_),
    .A2(_13469_),
    .B1(_13462_),
    .X(_13471_));
 sky130_fd_sc_hd__and3_1 _20193_ (.A(_13461_),
    .B(_13470_),
    .C(_13471_),
    .X(_13472_));
 sky130_fd_sc_hd__a21oi_1 _20194_ (.A1(_13470_),
    .A2(_13471_),
    .B1(_13461_),
    .Y(_13473_));
 sky130_fd_sc_hd__a211o_1 _20195_ (.A1(_13311_),
    .A2(_13313_),
    .B1(_13472_),
    .C1(_13473_),
    .X(_13474_));
 sky130_fd_sc_hd__o211ai_1 _20196_ (.A1(_13472_),
    .A2(_13473_),
    .B1(_13311_),
    .C1(_13313_),
    .Y(_13475_));
 sky130_fd_sc_hd__o211a_1 _20197_ (.A1(_13315_),
    .A2(_13317_),
    .B1(_13474_),
    .C1(_13475_),
    .X(_13476_));
 sky130_fd_sc_hd__a211oi_1 _20198_ (.A1(_13474_),
    .A2(_13475_),
    .B1(_13315_),
    .C1(_13317_),
    .Y(_13477_));
 sky130_fd_sc_hd__or4_2 _20199_ (.A(_13459_),
    .B(_13460_),
    .C(_13476_),
    .D(_13477_),
    .X(_13478_));
 sky130_fd_sc_hd__o22ai_2 _20200_ (.A1(_13459_),
    .A2(_13460_),
    .B1(_13476_),
    .B2(_13477_),
    .Y(_13479_));
 sky130_fd_sc_hd__o211ai_2 _20201_ (.A1(_13360_),
    .A2(_13362_),
    .B1(_13478_),
    .C1(_13479_),
    .Y(_13480_));
 sky130_fd_sc_hd__a211o_1 _20202_ (.A1(_13478_),
    .A2(_13479_),
    .B1(_13360_),
    .C1(_13362_),
    .X(_13481_));
 sky130_fd_sc_hd__o211a_1 _20203_ (.A1(_13319_),
    .A2(_13321_),
    .B1(_13480_),
    .C1(_13481_),
    .X(_13482_));
 sky130_fd_sc_hd__a211oi_1 _20204_ (.A1(_13480_),
    .A2(_13481_),
    .B1(_13319_),
    .C1(_13321_),
    .Y(_13483_));
 sky130_fd_sc_hd__clkbuf_4 _20205_ (.A(_12154_),
    .X(_13484_));
 sky130_fd_sc_hd__nand2_1 _20206_ (.A(_10893_),
    .B(_13484_),
    .Y(_13485_));
 sky130_fd_sc_hd__and4_1 _20207_ (.A(_11141_),
    .B(_11144_),
    .C(_12069_),
    .D(_12078_),
    .X(_13486_));
 sky130_fd_sc_hd__a22o_1 _20208_ (.A1(_11107_),
    .A2(_11958_),
    .B1(_12144_),
    .B2(_10956_),
    .X(_13487_));
 sky130_fd_sc_hd__and2b_1 _20209_ (.A_N(_13486_),
    .B(_13487_),
    .X(_13488_));
 sky130_fd_sc_hd__xnor2_2 _20210_ (.A(_13485_),
    .B(_13488_),
    .Y(_13489_));
 sky130_fd_sc_hd__nand2_1 _20211_ (.A(_11350_),
    .B(_11949_),
    .Y(_13490_));
 sky130_fd_sc_hd__nand4_2 _20212_ (.A(_11241_),
    .B(_11354_),
    .C(_11598_),
    .D(_12285_),
    .Y(_13491_));
 sky130_fd_sc_hd__a22o_1 _20213_ (.A1(_11458_),
    .A2(_11698_),
    .B1(_11707_),
    .B2(_11241_),
    .X(_13492_));
 sky130_fd_sc_hd__nand3b_1 _20214_ (.A_N(_13490_),
    .B(_13491_),
    .C(_13492_),
    .Y(_13493_));
 sky130_fd_sc_hd__a21bo_1 _20215_ (.A1(_13491_),
    .A2(_13492_),
    .B1_N(_13490_),
    .X(_13494_));
 sky130_fd_sc_hd__o21bai_1 _20216_ (.A1(_13335_),
    .A2(_13337_),
    .B1_N(_13336_),
    .Y(_13495_));
 sky130_fd_sc_hd__nand3_1 _20217_ (.A(_13493_),
    .B(_13494_),
    .C(_13495_),
    .Y(_13496_));
 sky130_fd_sc_hd__a21o_1 _20218_ (.A1(_13493_),
    .A2(_13494_),
    .B1(_13495_),
    .X(_13497_));
 sky130_fd_sc_hd__and3_1 _20219_ (.A(_13489_),
    .B(_13496_),
    .C(_13497_),
    .X(_13498_));
 sky130_fd_sc_hd__a21oi_1 _20220_ (.A1(_13496_),
    .A2(_13497_),
    .B1(_13489_),
    .Y(_13499_));
 sky130_fd_sc_hd__or2_1 _20221_ (.A(_13498_),
    .B(_13499_),
    .X(_13500_));
 sky130_fd_sc_hd__nand2_1 _20222_ (.A(_13347_),
    .B(_13349_),
    .Y(_13501_));
 sky130_fd_sc_hd__a31o_1 _20223_ (.A1(_11264_),
    .A2(_11770_),
    .A3(_13370_),
    .B1(_13369_),
    .X(_13502_));
 sky130_fd_sc_hd__nand2_1 _20224_ (.A(_11559_),
    .B(_11590_),
    .Y(_13503_));
 sky130_fd_sc_hd__nand4_2 _20225_ (.A(_11372_),
    .B(_11476_),
    .C(_11923_),
    .D(_11781_),
    .Y(_13504_));
 sky130_fd_sc_hd__a22o_1 _20226_ (.A1(_11476_),
    .A2(_11555_),
    .B1(_11658_),
    .B2(_11712_),
    .X(_13505_));
 sky130_fd_sc_hd__nand3b_1 _20227_ (.A_N(_13503_),
    .B(_13504_),
    .C(_13505_),
    .Y(_13506_));
 sky130_fd_sc_hd__a21bo_1 _20228_ (.A1(_13504_),
    .A2(_13505_),
    .B1_N(_13503_),
    .X(_13507_));
 sky130_fd_sc_hd__nand3_1 _20229_ (.A(_13502_),
    .B(_13506_),
    .C(_13507_),
    .Y(_13508_));
 sky130_fd_sc_hd__a21o_1 _20230_ (.A1(_13506_),
    .A2(_13507_),
    .B1(_13502_),
    .X(_13509_));
 sky130_fd_sc_hd__nand3_1 _20231_ (.A(_13501_),
    .B(_13508_),
    .C(_13509_),
    .Y(_13510_));
 sky130_fd_sc_hd__a21o_1 _20232_ (.A1(_13508_),
    .A2(_13509_),
    .B1(_13501_),
    .X(_13511_));
 sky130_fd_sc_hd__a21bo_1 _20233_ (.A1(_13345_),
    .A2(_13352_),
    .B1_N(_13351_),
    .X(_13512_));
 sky130_fd_sc_hd__and3_1 _20234_ (.A(_13510_),
    .B(_13511_),
    .C(_13512_),
    .X(_13513_));
 sky130_fd_sc_hd__a21oi_1 _20235_ (.A1(_13510_),
    .A2(_13511_),
    .B1(_13512_),
    .Y(_13514_));
 sky130_fd_sc_hd__nor3_2 _20236_ (.A(_13500_),
    .B(_13513_),
    .C(_13514_),
    .Y(_13515_));
 sky130_fd_sc_hd__o21a_1 _20237_ (.A1(_13513_),
    .A2(_13514_),
    .B1(_13500_),
    .X(_13516_));
 sky130_fd_sc_hd__a211o_1 _20238_ (.A1(_13385_),
    .A2(_13387_),
    .B1(_13515_),
    .C1(_13516_),
    .X(_13517_));
 sky130_fd_sc_hd__o211ai_1 _20239_ (.A1(_13515_),
    .A2(_13516_),
    .B1(_13385_),
    .C1(_13387_),
    .Y(_13518_));
 sky130_fd_sc_hd__o211a_1 _20240_ (.A1(_13356_),
    .A2(_13358_),
    .B1(_13517_),
    .C1(_13518_),
    .X(_13519_));
 sky130_fd_sc_hd__a211oi_1 _20241_ (.A1(_13517_),
    .A2(_13518_),
    .B1(_13356_),
    .C1(_13358_),
    .Y(_13520_));
 sky130_fd_sc_hd__a21bo_1 _20242_ (.A1(_13394_),
    .A2(_13401_),
    .B1_N(_13400_),
    .X(_13521_));
 sky130_fd_sc_hd__nand2_1 _20243_ (.A(_11172_),
    .B(_11895_),
    .Y(_13522_));
 sky130_fd_sc_hd__and4_1 _20244_ (.A(_11155_),
    .B(_11159_),
    .C(_12235_),
    .D(_12233_),
    .X(_13523_));
 sky130_fd_sc_hd__a22o_1 _20245_ (.A1(_11159_),
    .A2(_12235_),
    .B1(_12233_),
    .B2(_11155_),
    .X(_13524_));
 sky130_fd_sc_hd__and2b_1 _20246_ (.A_N(_13523_),
    .B(_13524_),
    .X(_13525_));
 sky130_fd_sc_hd__xnor2_2 _20247_ (.A(_13522_),
    .B(_13525_),
    .Y(_13526_));
 sky130_fd_sc_hd__nand2_1 _20248_ (.A(_10969_),
    .B(_12460_),
    .Y(_13527_));
 sky130_fd_sc_hd__and4_1 _20249_ (.A(_10909_),
    .B(_11174_),
    .C(_12327_),
    .D(_12600_),
    .X(_13528_));
 sky130_fd_sc_hd__a22oi_2 _20250_ (.A1(_10967_),
    .A2(_12322_),
    .B1(_13376_),
    .B2(_10852_),
    .Y(_13529_));
 sky130_fd_sc_hd__or3_1 _20251_ (.A(_13527_),
    .B(_13528_),
    .C(_13529_),
    .X(_13530_));
 sky130_fd_sc_hd__o21ai_1 _20252_ (.A1(_13528_),
    .A2(_13529_),
    .B1(_13527_),
    .Y(_13531_));
 sky130_fd_sc_hd__a21bo_1 _20253_ (.A1(_13373_),
    .A2(_13377_),
    .B1_N(_13375_),
    .X(_13532_));
 sky130_fd_sc_hd__nand3_1 _20254_ (.A(_13530_),
    .B(_13531_),
    .C(_13532_),
    .Y(_13533_));
 sky130_fd_sc_hd__a21o_1 _20255_ (.A1(_13530_),
    .A2(_13531_),
    .B1(_13532_),
    .X(_13534_));
 sky130_fd_sc_hd__nand3_1 _20256_ (.A(_13526_),
    .B(_13533_),
    .C(_13534_),
    .Y(_13535_));
 sky130_fd_sc_hd__a21o_1 _20257_ (.A1(_13533_),
    .A2(_13534_),
    .B1(_13526_),
    .X(_13536_));
 sky130_fd_sc_hd__and3_1 _20258_ (.A(_13521_),
    .B(_13535_),
    .C(_13536_),
    .X(_13537_));
 sky130_fd_sc_hd__a21oi_1 _20259_ (.A1(_13535_),
    .A2(_13536_),
    .B1(_13521_),
    .Y(_13538_));
 sky130_fd_sc_hd__a211oi_2 _20260_ (.A1(_13381_),
    .A2(_13383_),
    .B1(_13537_),
    .C1(_13538_),
    .Y(_13539_));
 sky130_fd_sc_hd__o211a_1 _20261_ (.A1(_13537_),
    .A2(_13538_),
    .B1(_13381_),
    .C1(_13383_),
    .X(_13540_));
 sky130_fd_sc_hd__clkbuf_2 _20262_ (.A(\genblk1.pcpi_mul.rs2[30] ),
    .X(_13541_));
 sky130_fd_sc_hd__and2_1 _20263_ (.A(_11113_),
    .B(_13541_),
    .X(_13542_));
 sky130_fd_sc_hd__nand2_1 _20264_ (.A(_10649_),
    .B(_13054_),
    .Y(_13543_));
 sky130_fd_sc_hd__and4_1 _20265_ (.A(_10786_),
    .B(_10754_),
    .C(\genblk1.pcpi_mul.rs2[28] ),
    .D(\genblk1.pcpi_mul.rs2[29] ),
    .X(_13544_));
 sky130_fd_sc_hd__clkbuf_2 _20266_ (.A(\genblk1.pcpi_mul.rs2[29] ),
    .X(_13545_));
 sky130_fd_sc_hd__a22oi_2 _20267_ (.A1(_11777_),
    .A2(_13227_),
    .B1(_13545_),
    .B2(_10705_),
    .Y(_13546_));
 sky130_fd_sc_hd__or3_1 _20268_ (.A(_13543_),
    .B(_13544_),
    .C(_13546_),
    .X(_13547_));
 sky130_fd_sc_hd__o21ai_1 _20269_ (.A1(_13544_),
    .A2(_13546_),
    .B1(_13543_),
    .Y(_13548_));
 sky130_fd_sc_hd__and3_1 _20270_ (.A(_13542_),
    .B(_13547_),
    .C(_13548_),
    .X(_13549_));
 sky130_fd_sc_hd__a21oi_1 _20271_ (.A1(_13547_),
    .A2(_13548_),
    .B1(_13542_),
    .Y(_13550_));
 sky130_fd_sc_hd__nor2_1 _20272_ (.A(_13549_),
    .B(_13550_),
    .Y(_13551_));
 sky130_fd_sc_hd__nand2_1 _20273_ (.A(_13396_),
    .B(_13398_),
    .Y(_13552_));
 sky130_fd_sc_hd__a31o_1 _20274_ (.A1(_11778_),
    .A2(_13054_),
    .A3(_13391_),
    .B1(_13390_),
    .X(_13553_));
 sky130_fd_sc_hd__nand2_1 _20275_ (.A(_10912_),
    .B(_12775_),
    .Y(_13554_));
 sky130_fd_sc_hd__buf_2 _20276_ (.A(_12770_),
    .X(_13555_));
 sky130_fd_sc_hd__clkbuf_2 _20277_ (.A(_12910_),
    .X(_13556_));
 sky130_fd_sc_hd__nand4_2 _20278_ (.A(_10742_),
    .B(_10697_),
    .C(_13555_),
    .D(_13556_),
    .Y(_13557_));
 sky130_fd_sc_hd__clkbuf_2 _20279_ (.A(_12909_),
    .X(_13558_));
 sky130_fd_sc_hd__a22o_1 _20280_ (.A1(_10746_),
    .A2(_13558_),
    .B1(_13556_),
    .B2(_10744_),
    .X(_13559_));
 sky130_fd_sc_hd__nand3b_1 _20281_ (.A_N(_13554_),
    .B(_13557_),
    .C(_13559_),
    .Y(_13560_));
 sky130_fd_sc_hd__a21bo_1 _20282_ (.A1(_13557_),
    .A2(_13559_),
    .B1_N(_13554_),
    .X(_13561_));
 sky130_fd_sc_hd__nand3_1 _20283_ (.A(_13553_),
    .B(_13560_),
    .C(_13561_),
    .Y(_13562_));
 sky130_fd_sc_hd__a21o_1 _20284_ (.A1(_13560_),
    .A2(_13561_),
    .B1(_13553_),
    .X(_13563_));
 sky130_fd_sc_hd__nand3_1 _20285_ (.A(_13552_),
    .B(_13562_),
    .C(_13563_),
    .Y(_13564_));
 sky130_fd_sc_hd__a21o_1 _20286_ (.A1(_13562_),
    .A2(_13563_),
    .B1(_13552_),
    .X(_13565_));
 sky130_fd_sc_hd__nand3_1 _20287_ (.A(_13551_),
    .B(_13564_),
    .C(_13565_),
    .Y(_13566_));
 sky130_fd_sc_hd__a21o_1 _20288_ (.A1(_13564_),
    .A2(_13565_),
    .B1(_13551_),
    .X(_13567_));
 sky130_fd_sc_hd__and3_1 _20289_ (.A(_13404_),
    .B(_13566_),
    .C(_13567_),
    .X(_13568_));
 sky130_fd_sc_hd__a21oi_1 _20290_ (.A1(_13566_),
    .A2(_13567_),
    .B1(_13404_),
    .Y(_13569_));
 sky130_fd_sc_hd__nor4_1 _20291_ (.A(_13539_),
    .B(_13540_),
    .C(_13568_),
    .D(_13569_),
    .Y(_13570_));
 sky130_fd_sc_hd__o22a_1 _20292_ (.A1(_13539_),
    .A2(_13540_),
    .B1(_13568_),
    .B2(_13569_),
    .X(_13571_));
 sky130_fd_sc_hd__a211oi_2 _20293_ (.A1(_13407_),
    .A2(_13409_),
    .B1(net361),
    .C1(_13571_),
    .Y(_13572_));
 sky130_fd_sc_hd__o211a_1 _20294_ (.A1(net361),
    .A2(_13571_),
    .B1(_13407_),
    .C1(_13409_),
    .X(_13573_));
 sky130_fd_sc_hd__nor4_1 _20295_ (.A(_13519_),
    .B(_13520_),
    .C(_13572_),
    .D(_13573_),
    .Y(_13574_));
 sky130_fd_sc_hd__o22a_1 _20296_ (.A1(_13519_),
    .A2(_13520_),
    .B1(_13572_),
    .B2(_13573_),
    .X(_13575_));
 sky130_fd_sc_hd__a211oi_2 _20297_ (.A1(_13411_),
    .A2(_13413_),
    .B1(net348),
    .C1(_13575_),
    .Y(_13576_));
 sky130_fd_sc_hd__o211a_1 _20298_ (.A1(net349),
    .A2(_13575_),
    .B1(_13411_),
    .C1(_13413_),
    .X(_13577_));
 sky130_fd_sc_hd__nor4_1 _20299_ (.A(_13482_),
    .B(_13483_),
    .C(_13576_),
    .D(_13577_),
    .Y(_13578_));
 sky130_fd_sc_hd__o22a_1 _20300_ (.A1(_13482_),
    .A2(_13483_),
    .B1(_13576_),
    .B2(_13577_),
    .X(_13579_));
 sky130_fd_sc_hd__a211oi_1 _20301_ (.A1(_13415_),
    .A2(_13417_),
    .B1(net340),
    .C1(_13579_),
    .Y(_13580_));
 sky130_fd_sc_hd__o211a_1 _20302_ (.A1(net340),
    .A2(_13579_),
    .B1(_13415_),
    .C1(_13417_),
    .X(_13581_));
 sky130_fd_sc_hd__or3_2 _20303_ (.A(_13436_),
    .B(_13580_),
    .C(_13581_),
    .X(_13582_));
 sky130_fd_sc_hd__o21ai_1 _20304_ (.A1(_13580_),
    .A2(_13581_),
    .B1(_13436_),
    .Y(_13583_));
 sky130_fd_sc_hd__o211a_1 _20305_ (.A1(_13419_),
    .A2(_13432_),
    .B1(_13582_),
    .C1(_13583_),
    .X(_13584_));
 sky130_fd_sc_hd__a211oi_1 _20306_ (.A1(_13582_),
    .A2(_13583_),
    .B1(_13419_),
    .C1(_13432_),
    .Y(_13585_));
 sky130_fd_sc_hd__or3_1 _20307_ (.A(_13269_),
    .B(_13584_),
    .C(_13585_),
    .X(_13586_));
 sky130_fd_sc_hd__o21ai_1 _20308_ (.A1(_13584_),
    .A2(_13585_),
    .B1(_13269_),
    .Y(_13587_));
 sky130_fd_sc_hd__nand2_2 _20309_ (.A(_13586_),
    .B(_13587_),
    .Y(_13588_));
 sky130_fd_sc_hd__and2b_1 _20310_ (.A_N(_13423_),
    .B(_13425_),
    .X(_13589_));
 sky130_fd_sc_hd__xor2_4 _20311_ (.A(_13588_),
    .B(_13589_),
    .X(_13590_));
 sky130_vsdinv _20312_ (.A(_13427_),
    .Y(_13591_));
 sky130_fd_sc_hd__a21o_1 _20313_ (.A1(_13430_),
    .A2(_13591_),
    .B1(_13428_),
    .X(_13592_));
 sky130_fd_sc_hd__o31ai_2 _20314_ (.A1(_13261_),
    .A2(_13265_),
    .A3(_13429_),
    .B1(_13592_),
    .Y(_13593_));
 sky130_fd_sc_hd__xor2_1 _20315_ (.A(_13590_),
    .B(_13593_),
    .X(_00076_));
 sky130_vsdinv _20316_ (.A(_13580_),
    .Y(_13594_));
 sky130_vsdinv _20317_ (.A(_13480_),
    .Y(_13595_));
 sky130_fd_sc_hd__nor2_1 _20318_ (.A(_13595_),
    .B(_13482_),
    .Y(_13596_));
 sky130_fd_sc_hd__nor2_1 _20319_ (.A(_13457_),
    .B(_13459_),
    .Y(_13597_));
 sky130_fd_sc_hd__xnor2_1 _20320_ (.A(_13596_),
    .B(_13597_),
    .Y(_13598_));
 sky130_vsdinv _20321_ (.A(_13478_),
    .Y(_13599_));
 sky130_fd_sc_hd__a211oi_2 _20322_ (.A1(_13385_),
    .A2(_13387_),
    .B1(_13515_),
    .C1(_13516_),
    .Y(_13600_));
 sky130_fd_sc_hd__or2_1 _20323_ (.A(_13280_),
    .B(_13442_),
    .X(_13601_));
 sky130_fd_sc_hd__a211o_1 _20324_ (.A1(_13282_),
    .A2(_13441_),
    .B1(_13443_),
    .C1(_13447_),
    .X(_13602_));
 sky130_fd_sc_hd__or2b_1 _20325_ (.A(_13454_),
    .B_N(_13453_),
    .X(_13603_));
 sky130_fd_sc_hd__nand2_1 _20326_ (.A(_13448_),
    .B(_13455_),
    .Y(_13604_));
 sky130_fd_sc_hd__clkbuf_2 _20327_ (.A(\genblk1.pcpi_mul.rs1[30] ),
    .X(_13605_));
 sky130_fd_sc_hd__clkbuf_2 _20328_ (.A(_13605_),
    .X(_13606_));
 sky130_fd_sc_hd__nand2_1 _20329_ (.A(_10627_),
    .B(_13606_),
    .Y(_13607_));
 sky130_fd_sc_hd__buf_2 _20330_ (.A(\genblk1.pcpi_mul.rs1[29] ),
    .X(_13608_));
 sky130_fd_sc_hd__clkbuf_2 _20331_ (.A(\genblk1.pcpi_mul.rs1[30] ),
    .X(_13609_));
 sky130_fd_sc_hd__and4_1 _20332_ (.A(_11044_),
    .B(_11041_),
    .C(_13608_),
    .D(_13609_),
    .X(_13610_));
 sky130_fd_sc_hd__a21oi_2 _20333_ (.A1(_13442_),
    .A2(_13607_),
    .B1(_13610_),
    .Y(_13611_));
 sky130_fd_sc_hd__buf_2 _20334_ (.A(_13281_),
    .X(_13612_));
 sky130_fd_sc_hd__nand2_2 _20335_ (.A(_10645_),
    .B(_13612_),
    .Y(_13613_));
 sky130_fd_sc_hd__xnor2_4 _20336_ (.A(_13611_),
    .B(_13613_),
    .Y(_13614_));
 sky130_fd_sc_hd__a22oi_2 _20337_ (.A1(_11061_),
    .A2(_12973_),
    .B1(_12980_),
    .B2(_11057_),
    .Y(_13615_));
 sky130_fd_sc_hd__and4_1 _20338_ (.A(_10671_),
    .B(_11711_),
    .C(_12973_),
    .D(\genblk1.pcpi_mul.rs1[27] ),
    .X(_13616_));
 sky130_fd_sc_hd__nor2_2 _20339_ (.A(_13615_),
    .B(_13616_),
    .Y(_13617_));
 sky130_fd_sc_hd__buf_2 _20340_ (.A(\genblk1.pcpi_mul.rs1[31] ),
    .X(_13618_));
 sky130_fd_sc_hd__nand2_2 _20341_ (.A(_11053_),
    .B(_13618_),
    .Y(_13619_));
 sky130_fd_sc_hd__xnor2_4 _20342_ (.A(_13617_),
    .B(_13619_),
    .Y(_13620_));
 sky130_fd_sc_hd__o21ba_1 _20343_ (.A1(_13449_),
    .A2(_13452_),
    .B1_N(_13450_),
    .X(_13621_));
 sky130_fd_sc_hd__xnor2_1 _20344_ (.A(_13620_),
    .B(_13621_),
    .Y(_13622_));
 sky130_fd_sc_hd__xnor2_1 _20345_ (.A(_13614_),
    .B(_13622_),
    .Y(_13623_));
 sky130_fd_sc_hd__a21oi_1 _20346_ (.A1(_13603_),
    .A2(_13604_),
    .B1(_13623_),
    .Y(_13624_));
 sky130_fd_sc_hd__and3_1 _20347_ (.A(_13603_),
    .B(_13604_),
    .C(_13623_),
    .X(_13625_));
 sky130_fd_sc_hd__a211oi_1 _20348_ (.A1(_13601_),
    .A2(_13602_),
    .B1(_13624_),
    .C1(_13625_),
    .Y(_13626_));
 sky130_fd_sc_hd__o211a_1 _20349_ (.A1(_13624_),
    .A2(_13625_),
    .B1(_13601_),
    .C1(_13602_),
    .X(_13627_));
 sky130_fd_sc_hd__nand3_1 _20350_ (.A(_13461_),
    .B(_13470_),
    .C(_13471_),
    .Y(_13628_));
 sky130_fd_sc_hd__a21bo_1 _20351_ (.A1(_13489_),
    .A2(_13497_),
    .B1_N(_13496_),
    .X(_13629_));
 sky130_fd_sc_hd__nand2_1 _20352_ (.A(_13465_),
    .B(_13467_),
    .Y(_13630_));
 sky130_fd_sc_hd__a31o_1 _20353_ (.A1(_10961_),
    .A2(_12274_),
    .A3(_13487_),
    .B1(_13486_),
    .X(_13631_));
 sky130_fd_sc_hd__buf_2 _20354_ (.A(_12700_),
    .X(_13632_));
 sky130_fd_sc_hd__a22o_1 _20355_ (.A1(_11196_),
    .A2(_12537_),
    .B1(_12688_),
    .B2(_11082_),
    .X(_13633_));
 sky130_fd_sc_hd__nand4_4 _20356_ (.A(_11298_),
    .B(_11086_),
    .C(_12538_),
    .D(_12690_),
    .Y(_13634_));
 sky130_fd_sc_hd__a22o_1 _20357_ (.A1(_11089_),
    .A2(_13632_),
    .B1(_13633_),
    .B2(_13634_),
    .X(_13635_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20358_ (.A(\genblk1.pcpi_mul.rs1[25] ),
    .X(_13636_));
 sky130_fd_sc_hd__clkbuf_4 _20359_ (.A(_13636_),
    .X(_13637_));
 sky130_fd_sc_hd__nand4_4 _20360_ (.A(_10737_),
    .B(_13637_),
    .C(_13633_),
    .D(_13634_),
    .Y(_13638_));
 sky130_fd_sc_hd__nand3_2 _20361_ (.A(_13631_),
    .B(_13635_),
    .C(_13638_),
    .Y(_13639_));
 sky130_fd_sc_hd__a21o_1 _20362_ (.A1(_13635_),
    .A2(_13638_),
    .B1(_13631_),
    .X(_13640_));
 sky130_fd_sc_hd__nand3_1 _20363_ (.A(_13630_),
    .B(_13639_),
    .C(_13640_),
    .Y(_13641_));
 sky130_fd_sc_hd__a21o_1 _20364_ (.A1(_13639_),
    .A2(_13640_),
    .B1(_13630_),
    .X(_13642_));
 sky130_fd_sc_hd__and3_1 _20365_ (.A(_13629_),
    .B(_13641_),
    .C(_13642_),
    .X(_13643_));
 sky130_fd_sc_hd__a21oi_1 _20366_ (.A1(_13641_),
    .A2(_13642_),
    .B1(_13629_),
    .Y(_13644_));
 sky130_fd_sc_hd__a211oi_2 _20367_ (.A1(_13468_),
    .A2(_13470_),
    .B1(_13643_),
    .C1(_13644_),
    .Y(_13645_));
 sky130_fd_sc_hd__o211a_1 _20368_ (.A1(_13643_),
    .A2(_13644_),
    .B1(_13468_),
    .C1(_13470_),
    .X(_13646_));
 sky130_fd_sc_hd__a211o_1 _20369_ (.A1(_13628_),
    .A2(_13474_),
    .B1(_13645_),
    .C1(_13646_),
    .X(_13647_));
 sky130_fd_sc_hd__o211ai_1 _20370_ (.A1(_13645_),
    .A2(_13646_),
    .B1(_13628_),
    .C1(_13474_),
    .Y(_13648_));
 sky130_fd_sc_hd__or4bb_1 _20371_ (.A(_13626_),
    .B(_13627_),
    .C_N(_13647_),
    .D_N(_13648_),
    .X(_13649_));
 sky130_fd_sc_hd__a2bb2o_1 _20372_ (.A1_N(_13626_),
    .A2_N(_13627_),
    .B1(_13647_),
    .B2(_13648_),
    .X(_13650_));
 sky130_fd_sc_hd__o211ai_2 _20373_ (.A1(_13600_),
    .A2(_13519_),
    .B1(_13649_),
    .C1(_13650_),
    .Y(_13651_));
 sky130_fd_sc_hd__a211o_1 _20374_ (.A1(_13649_),
    .A2(_13650_),
    .B1(_13600_),
    .C1(_13519_),
    .X(_13652_));
 sky130_fd_sc_hd__o211ai_2 _20375_ (.A1(_13476_),
    .A2(_13599_),
    .B1(_13651_),
    .C1(_13652_),
    .Y(_13653_));
 sky130_fd_sc_hd__a211o_1 _20376_ (.A1(_13651_),
    .A2(_13652_),
    .B1(_13476_),
    .C1(_13599_),
    .X(_13654_));
 sky130_vsdinv _20377_ (.A(_13572_),
    .Y(_13655_));
 sky130_fd_sc_hd__or4_1 _20378_ (.A(_13519_),
    .B(_13520_),
    .C(_13572_),
    .D(_13573_),
    .X(_13656_));
 sky130_vsdinv _20379_ (.A(_13513_),
    .Y(_13657_));
 sky130_vsdinv _20380_ (.A(_13515_),
    .Y(_13658_));
 sky130_fd_sc_hd__buf_2 _20381_ (.A(_12694_),
    .X(_13659_));
 sky130_fd_sc_hd__nand2_2 _20382_ (.A(_10894_),
    .B(_13659_),
    .Y(_13660_));
 sky130_fd_sc_hd__clkbuf_2 _20383_ (.A(_11142_),
    .X(_13661_));
 sky130_fd_sc_hd__clkbuf_2 _20384_ (.A(_11145_),
    .X(_13662_));
 sky130_fd_sc_hd__clkbuf_4 _20385_ (.A(_12144_),
    .X(_13663_));
 sky130_fd_sc_hd__and4_1 _20386_ (.A(_13661_),
    .B(_13662_),
    .C(_13663_),
    .D(_12543_),
    .X(_13664_));
 sky130_fd_sc_hd__buf_2 _20387_ (.A(_11108_),
    .X(_13665_));
 sky130_fd_sc_hd__buf_2 _20388_ (.A(_12147_),
    .X(_13666_));
 sky130_fd_sc_hd__buf_2 _20389_ (.A(_13666_),
    .X(_13667_));
 sky130_fd_sc_hd__clkbuf_4 _20390_ (.A(_12154_),
    .X(_13668_));
 sky130_fd_sc_hd__clkbuf_2 _20391_ (.A(_10963_),
    .X(_13669_));
 sky130_fd_sc_hd__buf_2 _20392_ (.A(_13669_),
    .X(_13670_));
 sky130_fd_sc_hd__a22oi_2 _20393_ (.A1(_13665_),
    .A2(_13667_),
    .B1(_13668_),
    .B2(_13670_),
    .Y(_13671_));
 sky130_fd_sc_hd__nor2_2 _20394_ (.A(_13664_),
    .B(_13671_),
    .Y(_13672_));
 sky130_fd_sc_hd__xnor2_4 _20395_ (.A(_13660_),
    .B(_13672_),
    .Y(_13673_));
 sky130_fd_sc_hd__buf_2 _20396_ (.A(_12067_),
    .X(_13674_));
 sky130_fd_sc_hd__nand2_2 _20397_ (.A(_11136_),
    .B(_13674_),
    .Y(_13675_));
 sky130_fd_sc_hd__clkbuf_2 _20398_ (.A(_11353_),
    .X(_13676_));
 sky130_fd_sc_hd__and4_1 _20399_ (.A(_11236_),
    .B(_13676_),
    .C(_11819_),
    .D(_11949_),
    .X(_13677_));
 sky130_fd_sc_hd__clkbuf_2 _20400_ (.A(_11354_),
    .X(_13678_));
 sky130_fd_sc_hd__buf_2 _20401_ (.A(_11946_),
    .X(_13679_));
 sky130_fd_sc_hd__clkbuf_2 _20402_ (.A(_11241_),
    .X(_13680_));
 sky130_fd_sc_hd__a22oi_2 _20403_ (.A1(_13678_),
    .A2(_11708_),
    .B1(_13679_),
    .B2(_13680_),
    .Y(_13681_));
 sky130_fd_sc_hd__nor2_2 _20404_ (.A(_13677_),
    .B(_13681_),
    .Y(_13682_));
 sky130_fd_sc_hd__xnor2_4 _20405_ (.A(_13675_),
    .B(_13682_),
    .Y(_13683_));
 sky130_fd_sc_hd__nand2_1 _20406_ (.A(_13491_),
    .B(_13493_),
    .Y(_13684_));
 sky130_fd_sc_hd__xor2_1 _20407_ (.A(_13683_),
    .B(_13684_),
    .X(_13685_));
 sky130_fd_sc_hd__xnor2_1 _20408_ (.A(_13673_),
    .B(_13685_),
    .Y(_13686_));
 sky130_fd_sc_hd__nand2_1 _20409_ (.A(_13504_),
    .B(_13506_),
    .Y(_13687_));
 sky130_fd_sc_hd__a31o_1 _20410_ (.A1(_11262_),
    .A2(_12591_),
    .A3(_13524_),
    .B1(_13523_),
    .X(_13688_));
 sky130_fd_sc_hd__clkbuf_4 _20411_ (.A(_12081_),
    .X(_13689_));
 sky130_fd_sc_hd__buf_2 _20412_ (.A(_13689_),
    .X(_13690_));
 sky130_fd_sc_hd__buf_2 _20413_ (.A(_11924_),
    .X(_13691_));
 sky130_fd_sc_hd__nand4_4 _20414_ (.A(_11834_),
    .B(_11590_),
    .C(_11663_),
    .D(_13691_),
    .Y(_13692_));
 sky130_fd_sc_hd__a22o_1 _20415_ (.A1(_11961_),
    .A2(_11923_),
    .B1(_11925_),
    .B2(_11380_),
    .X(_13693_));
 sky130_fd_sc_hd__nand4_4 _20416_ (.A(_11560_),
    .B(_13690_),
    .C(_13692_),
    .D(_13693_),
    .Y(_13694_));
 sky130_fd_sc_hd__clkbuf_2 _20417_ (.A(_11598_),
    .X(_13695_));
 sky130_fd_sc_hd__a22o_2 _20418_ (.A1(_11444_),
    .A2(_13695_),
    .B1(_13692_),
    .B2(_13693_),
    .X(_13696_));
 sky130_fd_sc_hd__nand3_2 _20419_ (.A(_13688_),
    .B(_13694_),
    .C(_13696_),
    .Y(_13697_));
 sky130_fd_sc_hd__a21o_1 _20420_ (.A1(_13694_),
    .A2(_13696_),
    .B1(_13688_),
    .X(_13698_));
 sky130_fd_sc_hd__nand3_1 _20421_ (.A(_13687_),
    .B(_13697_),
    .C(_13698_),
    .Y(_13699_));
 sky130_fd_sc_hd__a21o_1 _20422_ (.A1(_13697_),
    .A2(_13698_),
    .B1(_13687_),
    .X(_13700_));
 sky130_fd_sc_hd__a21bo_1 _20423_ (.A1(_13501_),
    .A2(_13509_),
    .B1_N(_13508_),
    .X(_13701_));
 sky130_fd_sc_hd__and3_1 _20424_ (.A(_13699_),
    .B(_13700_),
    .C(_13701_),
    .X(_13702_));
 sky130_fd_sc_hd__a21oi_1 _20425_ (.A1(_13699_),
    .A2(_13700_),
    .B1(_13701_),
    .Y(_13703_));
 sky130_fd_sc_hd__or3_1 _20426_ (.A(_13686_),
    .B(_13702_),
    .C(_13703_),
    .X(_13704_));
 sky130_fd_sc_hd__o21ai_1 _20427_ (.A1(_13702_),
    .A2(_13703_),
    .B1(_13686_),
    .Y(_13705_));
 sky130_fd_sc_hd__o211a_1 _20428_ (.A1(_13537_),
    .A2(_13539_),
    .B1(_13704_),
    .C1(_13705_),
    .X(_13706_));
 sky130_fd_sc_hd__a211oi_1 _20429_ (.A1(_13704_),
    .A2(_13705_),
    .B1(_13537_),
    .C1(_13539_),
    .Y(_13707_));
 sky130_fd_sc_hd__a211oi_2 _20430_ (.A1(_13657_),
    .A2(_13658_),
    .B1(_13706_),
    .C1(_13707_),
    .Y(_13708_));
 sky130_fd_sc_hd__o211a_1 _20431_ (.A1(_13706_),
    .A2(_13707_),
    .B1(_13657_),
    .C1(_13658_),
    .X(_13709_));
 sky130_fd_sc_hd__a21bo_1 _20432_ (.A1(_13552_),
    .A2(_13563_),
    .B1_N(_13562_),
    .X(_13710_));
 sky130_fd_sc_hd__buf_4 _20433_ (.A(_11895_),
    .X(_13711_));
 sky130_fd_sc_hd__nand2_1 _20434_ (.A(_11369_),
    .B(_13711_),
    .Y(_13712_));
 sky130_fd_sc_hd__buf_2 _20435_ (.A(_12235_),
    .X(_13713_));
 sky130_fd_sc_hd__and4_1 _20436_ (.A(_11728_),
    .B(_11265_),
    .C(_13713_),
    .D(_12023_),
    .X(_13714_));
 sky130_fd_sc_hd__buf_2 _20437_ (.A(_12233_),
    .X(_13715_));
 sky130_fd_sc_hd__clkbuf_4 _20438_ (.A(_13715_),
    .X(_13716_));
 sky130_fd_sc_hd__a22oi_4 _20439_ (.A1(_11172_),
    .A2(_11891_),
    .B1(_13716_),
    .B2(_11068_),
    .Y(_13717_));
 sky130_fd_sc_hd__nor2_1 _20440_ (.A(_13714_),
    .B(_13717_),
    .Y(_13718_));
 sky130_fd_sc_hd__xnor2_1 _20441_ (.A(_13712_),
    .B(_13718_),
    .Y(_13719_));
 sky130_fd_sc_hd__clkbuf_4 _20442_ (.A(_12226_),
    .X(_13720_));
 sky130_fd_sc_hd__clkbuf_4 _20443_ (.A(_13374_),
    .X(_13721_));
 sky130_fd_sc_hd__nand4_4 _20444_ (.A(_11049_),
    .B(_11042_),
    .C(_12329_),
    .D(_13721_),
    .Y(_13722_));
 sky130_fd_sc_hd__buf_2 _20445_ (.A(_12600_),
    .X(_13723_));
 sky130_fd_sc_hd__a22o_1 _20446_ (.A1(_11280_),
    .A2(_12323_),
    .B1(_13723_),
    .B2(_11177_),
    .X(_13724_));
 sky130_fd_sc_hd__nand4_2 _20447_ (.A(_11157_),
    .B(_13720_),
    .C(_13722_),
    .D(_13724_),
    .Y(_13725_));
 sky130_fd_sc_hd__a22o_1 _20448_ (.A1(_11270_),
    .A2(_12227_),
    .B1(_13722_),
    .B2(_13724_),
    .X(_13726_));
 sky130_fd_sc_hd__o21bai_1 _20449_ (.A1(_13527_),
    .A2(_13529_),
    .B1_N(_13528_),
    .Y(_13727_));
 sky130_fd_sc_hd__nand3_1 _20450_ (.A(_13725_),
    .B(_13726_),
    .C(_13727_),
    .Y(_13728_));
 sky130_fd_sc_hd__a21o_1 _20451_ (.A1(_13725_),
    .A2(_13726_),
    .B1(_13727_),
    .X(_13729_));
 sky130_fd_sc_hd__nand3_1 _20452_ (.A(_13719_),
    .B(_13728_),
    .C(_13729_),
    .Y(_13730_));
 sky130_fd_sc_hd__a21o_1 _20453_ (.A1(_13728_),
    .A2(_13729_),
    .B1(_13719_),
    .X(_13731_));
 sky130_fd_sc_hd__and3_1 _20454_ (.A(_13710_),
    .B(_13730_),
    .C(_13731_),
    .X(_13732_));
 sky130_fd_sc_hd__a21oi_1 _20455_ (.A1(_13730_),
    .A2(_13731_),
    .B1(_13710_),
    .Y(_13733_));
 sky130_fd_sc_hd__a211o_1 _20456_ (.A1(_13533_),
    .A2(_13535_),
    .B1(_13732_),
    .C1(_13733_),
    .X(_13734_));
 sky130_fd_sc_hd__o211ai_1 _20457_ (.A1(_13732_),
    .A2(_13733_),
    .B1(_13533_),
    .C1(_13535_),
    .Y(_13735_));
 sky130_fd_sc_hd__nand2_1 _20458_ (.A(_13557_),
    .B(_13560_),
    .Y(_13736_));
 sky130_fd_sc_hd__o21bai_1 _20459_ (.A1(_13543_),
    .A2(_13546_),
    .B1_N(_13544_),
    .Y(_13737_));
 sky130_fd_sc_hd__clkbuf_4 _20460_ (.A(_12584_),
    .X(_13738_));
 sky130_fd_sc_hd__clkbuf_4 _20461_ (.A(_13555_),
    .X(_13739_));
 sky130_fd_sc_hd__clkbuf_2 _20462_ (.A(\genblk1.pcpi_mul.rs2[26] ),
    .X(_13740_));
 sky130_fd_sc_hd__clkbuf_4 _20463_ (.A(_13740_),
    .X(_13741_));
 sky130_fd_sc_hd__nand4_2 _20464_ (.A(_11193_),
    .B(_11091_),
    .C(_13739_),
    .D(_13741_),
    .Y(_13742_));
 sky130_fd_sc_hd__clkbuf_4 _20465_ (.A(_13060_),
    .X(_13743_));
 sky130_fd_sc_hd__clkbuf_4 _20466_ (.A(_13740_),
    .X(_13744_));
 sky130_fd_sc_hd__a22o_1 _20467_ (.A1(_11302_),
    .A2(_13743_),
    .B1(_13744_),
    .B2(_10855_),
    .X(_13745_));
 sky130_fd_sc_hd__nand4_2 _20468_ (.A(_11297_),
    .B(_13738_),
    .C(_13742_),
    .D(_13745_),
    .Y(_13746_));
 sky130_fd_sc_hd__a22o_1 _20469_ (.A1(_11297_),
    .A2(_13738_),
    .B1(_13742_),
    .B2(_13745_),
    .X(_13747_));
 sky130_fd_sc_hd__nand3_2 _20470_ (.A(_13737_),
    .B(_13746_),
    .C(_13747_),
    .Y(_13748_));
 sky130_fd_sc_hd__a21o_1 _20471_ (.A1(_13746_),
    .A2(_13747_),
    .B1(_13737_),
    .X(_13749_));
 sky130_fd_sc_hd__nand3_1 _20472_ (.A(_13736_),
    .B(_13748_),
    .C(_13749_),
    .Y(_13750_));
 sky130_fd_sc_hd__a21o_1 _20473_ (.A1(_13748_),
    .A2(_13749_),
    .B1(_13736_),
    .X(_13751_));
 sky130_fd_sc_hd__clkbuf_2 _20474_ (.A(\genblk1.pcpi_mul.rs2[30] ),
    .X(_13752_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20475_ (.A(\genblk1.pcpi_mul.rs2[31] ),
    .X(_13753_));
 sky130_fd_sc_hd__clkbuf_4 _20476_ (.A(_13753_),
    .X(_13754_));
 sky130_fd_sc_hd__a22oi_1 _20477_ (.A1(_10636_),
    .A2(_13752_),
    .B1(_13754_),
    .B2(_10589_),
    .Y(_13755_));
 sky130_fd_sc_hd__clkbuf_2 _20478_ (.A(\genblk1.pcpi_mul.rs2[31] ),
    .X(_13756_));
 sky130_fd_sc_hd__buf_2 _20479_ (.A(_13756_),
    .X(_13757_));
 sky130_fd_sc_hd__and4_2 _20480_ (.A(_11113_),
    .B(_10638_),
    .C(_13541_),
    .D(_13757_),
    .X(_13758_));
 sky130_fd_sc_hd__nor2_1 _20481_ (.A(_13755_),
    .B(_13758_),
    .Y(_13759_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20482_ (.A(\genblk1.pcpi_mul.rs2[28] ),
    .X(_13760_));
 sky130_fd_sc_hd__clkbuf_2 _20483_ (.A(_13760_),
    .X(_13761_));
 sky130_fd_sc_hd__buf_2 _20484_ (.A(_13545_),
    .X(_13762_));
 sky130_fd_sc_hd__nand4_2 _20485_ (.A(_10608_),
    .B(_10676_),
    .C(_13761_),
    .D(_13762_),
    .Y(_13763_));
 sky130_fd_sc_hd__clkbuf_2 _20486_ (.A(_13227_),
    .X(_13764_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20487_ (.A(\genblk1.pcpi_mul.rs2[29] ),
    .X(_13765_));
 sky130_fd_sc_hd__a22o_1 _20488_ (.A1(_10650_),
    .A2(_13764_),
    .B1(_13765_),
    .B2(_11778_),
    .X(_13766_));
 sky130_fd_sc_hd__nand4_2 _20489_ (.A(_10667_),
    .B(_13056_),
    .C(_13763_),
    .D(_13766_),
    .Y(_13767_));
 sky130_fd_sc_hd__a22o_1 _20490_ (.A1(_11245_),
    .A2(_13226_),
    .B1(_13763_),
    .B2(_13766_),
    .X(_13768_));
 sky130_fd_sc_hd__nand3_4 _20491_ (.A(_13759_),
    .B(_13767_),
    .C(_13768_),
    .Y(_13769_));
 sky130_fd_sc_hd__a21o_1 _20492_ (.A1(_13767_),
    .A2(_13768_),
    .B1(_13759_),
    .X(_13770_));
 sky130_fd_sc_hd__nand3_1 _20493_ (.A(_13549_),
    .B(_13769_),
    .C(_13770_),
    .Y(_13771_));
 sky130_fd_sc_hd__a21o_1 _20494_ (.A1(_13769_),
    .A2(_13770_),
    .B1(_13549_),
    .X(_13772_));
 sky130_fd_sc_hd__nand4_1 _20495_ (.A(_13750_),
    .B(_13751_),
    .C(_13771_),
    .D(_13772_),
    .Y(_13773_));
 sky130_fd_sc_hd__a22o_1 _20496_ (.A1(_13750_),
    .A2(_13751_),
    .B1(_13771_),
    .B2(_13772_),
    .X(_13774_));
 sky130_fd_sc_hd__nand3b_1 _20497_ (.A_N(_13566_),
    .B(_13773_),
    .C(_13774_),
    .Y(_13775_));
 sky130_fd_sc_hd__a21bo_1 _20498_ (.A1(_13773_),
    .A2(_13774_),
    .B1_N(_13566_),
    .X(_13776_));
 sky130_fd_sc_hd__nand4_1 _20499_ (.A(_13734_),
    .B(_13735_),
    .C(_13775_),
    .D(_13776_),
    .Y(_13777_));
 sky130_fd_sc_hd__a22o_1 _20500_ (.A1(_13734_),
    .A2(_13735_),
    .B1(_13775_),
    .B2(_13776_),
    .X(_13778_));
 sky130_fd_sc_hd__o211a_1 _20501_ (.A1(_13568_),
    .A2(net418),
    .B1(_13777_),
    .C1(_13778_),
    .X(_13779_));
 sky130_fd_sc_hd__a211oi_1 _20502_ (.A1(_13777_),
    .A2(_13778_),
    .B1(_13568_),
    .C1(net418),
    .Y(_13780_));
 sky130_fd_sc_hd__nor4_2 _20503_ (.A(_13708_),
    .B(_13709_),
    .C(_13779_),
    .D(_13780_),
    .Y(_13781_));
 sky130_fd_sc_hd__o22a_1 _20504_ (.A1(_13708_),
    .A2(_13709_),
    .B1(_13779_),
    .B2(_13780_),
    .X(_13782_));
 sky130_fd_sc_hd__a211o_1 _20505_ (.A1(_13655_),
    .A2(_13656_),
    .B1(_13781_),
    .C1(_13782_),
    .X(_13783_));
 sky130_fd_sc_hd__o211ai_2 _20506_ (.A1(_13781_),
    .A2(_13782_),
    .B1(_13655_),
    .C1(_13656_),
    .Y(_13784_));
 sky130_fd_sc_hd__nand4_2 _20507_ (.A(_13653_),
    .B(_13654_),
    .C(_13783_),
    .D(_13784_),
    .Y(_13785_));
 sky130_fd_sc_hd__a22o_1 _20508_ (.A1(_13653_),
    .A2(_13654_),
    .B1(_13783_),
    .B2(_13784_),
    .X(_13786_));
 sky130_fd_sc_hd__o211a_1 _20509_ (.A1(_13576_),
    .A2(net415),
    .B1(_13785_),
    .C1(_13786_),
    .X(_13787_));
 sky130_fd_sc_hd__a211oi_1 _20510_ (.A1(_13785_),
    .A2(_13786_),
    .B1(_13576_),
    .C1(net415),
    .Y(_13788_));
 sky130_fd_sc_hd__nor3_2 _20511_ (.A(_13598_),
    .B(_13787_),
    .C(_13788_),
    .Y(_13789_));
 sky130_fd_sc_hd__o21a_1 _20512_ (.A1(_13787_),
    .A2(_13788_),
    .B1(_13598_),
    .X(_13790_));
 sky130_fd_sc_hd__a211oi_2 _20513_ (.A1(_13594_),
    .A2(_13582_),
    .B1(_13789_),
    .C1(_13790_),
    .Y(_13791_));
 sky130_fd_sc_hd__o211a_1 _20514_ (.A1(_13789_),
    .A2(_13790_),
    .B1(_13594_),
    .C1(_13582_),
    .X(_13792_));
 sky130_fd_sc_hd__nor3_1 _20515_ (.A(_13434_),
    .B(_13791_),
    .C(_13792_),
    .Y(_13793_));
 sky130_fd_sc_hd__o21a_1 _20516_ (.A1(_13791_),
    .A2(_13792_),
    .B1(_13434_),
    .X(_13794_));
 sky130_vsdinv _20517_ (.A(_13584_),
    .Y(_13795_));
 sky130_fd_sc_hd__o211a_1 _20518_ (.A1(net335),
    .A2(_13794_),
    .B1(_13795_),
    .C1(_13586_),
    .X(_13796_));
 sky130_fd_sc_hd__a211o_1 _20519_ (.A1(_13795_),
    .A2(_13586_),
    .B1(net335),
    .C1(_13794_),
    .X(_13797_));
 sky130_fd_sc_hd__nor2b_2 _20520_ (.A(_13796_),
    .B_N(_13797_),
    .Y(_13798_));
 sky130_fd_sc_hd__or2_2 _20521_ (.A(_13588_),
    .B(_13589_),
    .X(_13799_));
 sky130_fd_sc_hd__a21bo_1 _20522_ (.A1(_13590_),
    .A2(_13593_),
    .B1_N(_13799_),
    .X(_13800_));
 sky130_fd_sc_hd__xor2_1 _20523_ (.A(_13798_),
    .B(_13800_),
    .X(_00077_));
 sky130_fd_sc_hd__nor2_2 _20524_ (.A(_13596_),
    .B(_13597_),
    .Y(_13801_));
 sky130_fd_sc_hd__buf_1 _20525_ (.A(\genblk1.pcpi_mul.rs2[32] ),
    .X(_13802_));
 sky130_fd_sc_hd__buf_2 _20526_ (.A(_13802_),
    .X(_13803_));
 sky130_fd_sc_hd__clkbuf_2 _20527_ (.A(_13803_),
    .X(_13804_));
 sky130_fd_sc_hd__buf_4 _20528_ (.A(_13804_),
    .X(_13805_));
 sky130_fd_sc_hd__nor2_1 _20529_ (.A(_13624_),
    .B(_13626_),
    .Y(_13806_));
 sky130_fd_sc_hd__a21oi_1 _20530_ (.A1(_13651_),
    .A2(_13653_),
    .B1(_13806_),
    .Y(_13807_));
 sky130_fd_sc_hd__and3_1 _20531_ (.A(_13651_),
    .B(_13653_),
    .C(_13806_),
    .X(_13808_));
 sky130_fd_sc_hd__nor2_1 _20532_ (.A(_13807_),
    .B(_13808_),
    .Y(_13809_));
 sky130_fd_sc_hd__xnor2_1 _20533_ (.A(_13805_),
    .B(_13809_),
    .Y(_13810_));
 sky130_fd_sc_hd__nand2_1 _20534_ (.A(_13647_),
    .B(_13649_),
    .Y(_13811_));
 sky130_fd_sc_hd__or2_1 _20535_ (.A(_13706_),
    .B(_13708_),
    .X(_13812_));
 sky130_fd_sc_hd__clkbuf_2 _20536_ (.A(\genblk1.pcpi_mul.rs1[29] ),
    .X(_13813_));
 sky130_fd_sc_hd__buf_2 _20537_ (.A(_13813_),
    .X(_13814_));
 sky130_fd_sc_hd__clkbuf_4 _20538_ (.A(_13814_),
    .X(_13815_));
 sky130_fd_sc_hd__clkbuf_4 _20539_ (.A(_13815_),
    .X(_13816_));
 sky130_fd_sc_hd__buf_2 _20540_ (.A(_13606_),
    .X(_13817_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20541_ (.A(_13817_),
    .X(_13818_));
 sky130_fd_sc_hd__clkbuf_4 _20542_ (.A(_13818_),
    .X(_13819_));
 sky130_fd_sc_hd__nand4_4 _20543_ (.A(_10602_),
    .B(_10613_),
    .C(_13816_),
    .D(_13819_),
    .Y(_13820_));
 sky130_fd_sc_hd__a211o_2 _20544_ (.A1(_13442_),
    .A2(_13607_),
    .B1(_13610_),
    .C1(_13613_),
    .X(_13821_));
 sky130_fd_sc_hd__or2b_1 _20545_ (.A(_13621_),
    .B_N(_13620_),
    .X(_13822_));
 sky130_fd_sc_hd__nand2_1 _20546_ (.A(_13614_),
    .B(_13622_),
    .Y(_13823_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20547_ (.A(_13608_),
    .X(_13824_));
 sky130_fd_sc_hd__buf_2 _20548_ (.A(_13824_),
    .X(_13825_));
 sky130_fd_sc_hd__clkbuf_2 _20549_ (.A(_13609_),
    .X(_13826_));
 sky130_fd_sc_hd__buf_2 _20550_ (.A(_13618_),
    .X(_13827_));
 sky130_fd_sc_hd__a22o_1 _20551_ (.A1(_10613_),
    .A2(_13826_),
    .B1(_13827_),
    .B2(_10601_),
    .X(_13828_));
 sky130_fd_sc_hd__clkbuf_4 _20552_ (.A(_13606_),
    .X(_13829_));
 sky130_fd_sc_hd__clkbuf_2 _20553_ (.A(\genblk1.pcpi_mul.rs1[31] ),
    .X(_13830_));
 sky130_fd_sc_hd__clkbuf_4 _20554_ (.A(_13830_),
    .X(_13831_));
 sky130_fd_sc_hd__nand4_4 _20555_ (.A(_10601_),
    .B(_10613_),
    .C(_13829_),
    .D(_13831_),
    .Y(_13832_));
 sky130_fd_sc_hd__a22o_1 _20556_ (.A1(_10680_),
    .A2(_13825_),
    .B1(_13828_),
    .B2(_13832_),
    .X(_13833_));
 sky130_fd_sc_hd__nand4_2 _20557_ (.A(_10680_),
    .B(_13815_),
    .C(_13828_),
    .D(_13832_),
    .Y(_13834_));
 sky130_fd_sc_hd__and2_1 _20558_ (.A(_13833_),
    .B(_13834_),
    .X(_13835_));
 sky130_fd_sc_hd__clkbuf_2 _20559_ (.A(_13128_),
    .X(_13836_));
 sky130_fd_sc_hd__a22oi_1 _20560_ (.A1(_11385_),
    .A2(_13446_),
    .B1(_13836_),
    .B2(_11387_),
    .Y(_13837_));
 sky130_fd_sc_hd__clkbuf_2 _20561_ (.A(_12980_),
    .X(_13838_));
 sky130_fd_sc_hd__clkbuf_2 _20562_ (.A(_13128_),
    .X(_13839_));
 sky130_fd_sc_hd__and4_1 _20563_ (.A(_10672_),
    .B(_11282_),
    .C(_13838_),
    .D(_13839_),
    .X(_13840_));
 sky130_fd_sc_hd__nor2_1 _20564_ (.A(_13837_),
    .B(_13840_),
    .Y(_13841_));
 sky130_fd_sc_hd__buf_2 _20565_ (.A(\genblk1.pcpi_mul.rs1[32] ),
    .X(_13842_));
 sky130_fd_sc_hd__nand2_2 _20566_ (.A(_11053_),
    .B(_13842_),
    .Y(_13843_));
 sky130_fd_sc_hd__xnor2_1 _20567_ (.A(_13841_),
    .B(_13843_),
    .Y(_13844_));
 sky130_fd_sc_hd__o21ba_2 _20568_ (.A1(_13615_),
    .A2(_13619_),
    .B1_N(_13616_),
    .X(_13845_));
 sky130_fd_sc_hd__xnor2_1 _20569_ (.A(_13844_),
    .B(_13845_),
    .Y(_13846_));
 sky130_fd_sc_hd__and2_1 _20570_ (.A(_13835_),
    .B(_13846_),
    .X(_13847_));
 sky130_fd_sc_hd__nor2_1 _20571_ (.A(_13835_),
    .B(_13846_),
    .Y(_13848_));
 sky130_fd_sc_hd__or2_4 _20572_ (.A(_13847_),
    .B(_13848_),
    .X(_13849_));
 sky130_fd_sc_hd__a21oi_2 _20573_ (.A1(_13822_),
    .A2(_13823_),
    .B1(_13849_),
    .Y(_13850_));
 sky130_fd_sc_hd__and3_1 _20574_ (.A(_13822_),
    .B(_13823_),
    .C(_13849_),
    .X(_13851_));
 sky130_fd_sc_hd__a211oi_2 _20575_ (.A1(_13820_),
    .A2(_13821_),
    .B1(_13850_),
    .C1(_13851_),
    .Y(_13852_));
 sky130_fd_sc_hd__o211a_1 _20576_ (.A1(_13850_),
    .A2(_13851_),
    .B1(_13820_),
    .C1(_13821_),
    .X(_13853_));
 sky130_fd_sc_hd__and2_1 _20577_ (.A(_13683_),
    .B(_13684_),
    .X(_13854_));
 sky130_fd_sc_hd__and2_1 _20578_ (.A(_13673_),
    .B(_13685_),
    .X(_13855_));
 sky130_fd_sc_hd__nand2_2 _20579_ (.A(_13634_),
    .B(_13638_),
    .Y(_13856_));
 sky130_fd_sc_hd__o21ba_2 _20580_ (.A1(_13660_),
    .A2(_13671_),
    .B1_N(_13664_),
    .X(_13857_));
 sky130_fd_sc_hd__buf_4 _20581_ (.A(_11086_),
    .X(_13858_));
 sky130_fd_sc_hd__clkbuf_2 _20582_ (.A(_12688_),
    .X(_13859_));
 sky130_fd_sc_hd__buf_2 _20583_ (.A(_13859_),
    .X(_13860_));
 sky130_fd_sc_hd__buf_2 _20584_ (.A(_13632_),
    .X(_13861_));
 sky130_fd_sc_hd__a22oi_2 _20585_ (.A1(_13858_),
    .A2(_13860_),
    .B1(_13861_),
    .B2(_10784_),
    .Y(_13862_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20586_ (.A(_11084_),
    .X(_13863_));
 sky130_fd_sc_hd__buf_2 _20587_ (.A(_13632_),
    .X(_13864_));
 sky130_fd_sc_hd__and4_1 _20588_ (.A(_13863_),
    .B(_13858_),
    .C(_12977_),
    .D(_13864_),
    .X(_13865_));
 sky130_fd_sc_hd__nor2_2 _20589_ (.A(_13862_),
    .B(_13865_),
    .Y(_13866_));
 sky130_fd_sc_hd__clkbuf_2 _20590_ (.A(\genblk1.pcpi_mul.rs1[26] ),
    .X(_13867_));
 sky130_fd_sc_hd__clkbuf_2 _20591_ (.A(_13867_),
    .X(_13868_));
 sky130_fd_sc_hd__buf_2 _20592_ (.A(_13868_),
    .X(_13869_));
 sky130_fd_sc_hd__nand2_2 _20593_ (.A(_10738_),
    .B(_13869_),
    .Y(_13870_));
 sky130_fd_sc_hd__xnor2_4 _20594_ (.A(_13866_),
    .B(_13870_),
    .Y(_13871_));
 sky130_fd_sc_hd__xnor2_4 _20595_ (.A(_13857_),
    .B(_13871_),
    .Y(_13872_));
 sky130_fd_sc_hd__xor2_2 _20596_ (.A(_13856_),
    .B(_13872_),
    .X(_13873_));
 sky130_fd_sc_hd__o21a_1 _20597_ (.A1(_13854_),
    .A2(_13855_),
    .B1(_13873_),
    .X(_13874_));
 sky130_fd_sc_hd__nor3_1 _20598_ (.A(_13854_),
    .B(_13855_),
    .C(_13873_),
    .Y(_13875_));
 sky130_fd_sc_hd__a211o_1 _20599_ (.A1(_13639_),
    .A2(_13641_),
    .B1(_13874_),
    .C1(_13875_),
    .X(_13876_));
 sky130_fd_sc_hd__o211ai_1 _20600_ (.A1(_13874_),
    .A2(_13875_),
    .B1(_13639_),
    .C1(_13641_),
    .Y(_13877_));
 sky130_fd_sc_hd__o211a_1 _20601_ (.A1(_13643_),
    .A2(_13645_),
    .B1(_13876_),
    .C1(_13877_),
    .X(_13878_));
 sky130_fd_sc_hd__a211oi_1 _20602_ (.A1(_13876_),
    .A2(_13877_),
    .B1(_13643_),
    .C1(_13645_),
    .Y(_13879_));
 sky130_fd_sc_hd__nor4_1 _20603_ (.A(_13852_),
    .B(_13853_),
    .C(_13878_),
    .D(_13879_),
    .Y(_13880_));
 sky130_fd_sc_hd__o22a_1 _20604_ (.A1(_13852_),
    .A2(_13853_),
    .B1(_13878_),
    .B2(_13879_),
    .X(_13881_));
 sky130_fd_sc_hd__nor2_1 _20605_ (.A(_13880_),
    .B(_13881_),
    .Y(_13882_));
 sky130_fd_sc_hd__xnor2_1 _20606_ (.A(_13812_),
    .B(_13882_),
    .Y(_13883_));
 sky130_fd_sc_hd__xnor2_2 _20607_ (.A(_13811_),
    .B(_13883_),
    .Y(_13884_));
 sky130_fd_sc_hd__and2b_1 _20608_ (.A_N(_13702_),
    .B(_13704_),
    .X(_13885_));
 sky130_fd_sc_hd__nand3_1 _20609_ (.A(_13710_),
    .B(_13730_),
    .C(_13731_),
    .Y(_13886_));
 sky130_fd_sc_hd__clkbuf_2 _20610_ (.A(_12416_),
    .X(_13887_));
 sky130_fd_sc_hd__buf_2 _20611_ (.A(_13887_),
    .X(_13888_));
 sky130_fd_sc_hd__nand2_1 _20612_ (.A(_10894_),
    .B(_13888_),
    .Y(_13889_));
 sky130_fd_sc_hd__buf_2 _20613_ (.A(_12983_),
    .X(_13890_));
 sky130_fd_sc_hd__buf_2 _20614_ (.A(_13890_),
    .X(_13891_));
 sky130_fd_sc_hd__and4_1 _20615_ (.A(_13670_),
    .B(_13665_),
    .C(_13668_),
    .D(_13891_),
    .X(_13892_));
 sky130_fd_sc_hd__buf_2 _20616_ (.A(_13484_),
    .X(_13893_));
 sky130_fd_sc_hd__a22oi_4 _20617_ (.A1(_11109_),
    .A2(_13893_),
    .B1(_13659_),
    .B2(_10958_),
    .Y(_13894_));
 sky130_fd_sc_hd__nor2_1 _20618_ (.A(_13892_),
    .B(_13894_),
    .Y(_13895_));
 sky130_fd_sc_hd__xnor2_1 _20619_ (.A(_13889_),
    .B(_13895_),
    .Y(_13896_));
 sky130_fd_sc_hd__clkbuf_2 _20620_ (.A(_11135_),
    .X(_13897_));
 sky130_fd_sc_hd__nand2_1 _20621_ (.A(_13897_),
    .B(_13667_),
    .Y(_13898_));
 sky130_fd_sc_hd__clkbuf_2 _20622_ (.A(_11236_),
    .X(_13899_));
 sky130_fd_sc_hd__clkbuf_2 _20623_ (.A(_13676_),
    .X(_13900_));
 sky130_fd_sc_hd__buf_2 _20624_ (.A(_13305_),
    .X(_13901_));
 sky130_fd_sc_hd__and4_1 _20625_ (.A(_13899_),
    .B(_13900_),
    .C(_11831_),
    .D(_13901_),
    .X(_13902_));
 sky130_fd_sc_hd__buf_2 _20626_ (.A(_13676_),
    .X(_13903_));
 sky130_fd_sc_hd__buf_2 _20627_ (.A(_13679_),
    .X(_13904_));
 sky130_fd_sc_hd__a22oi_2 _20628_ (.A1(_13903_),
    .A2(_13904_),
    .B1(_13674_),
    .B2(_11237_),
    .Y(_13905_));
 sky130_fd_sc_hd__nor2_1 _20629_ (.A(_13902_),
    .B(_13905_),
    .Y(_13906_));
 sky130_fd_sc_hd__xnor2_1 _20630_ (.A(_13898_),
    .B(_13906_),
    .Y(_13907_));
 sky130_fd_sc_hd__o21ba_1 _20631_ (.A1(_13675_),
    .A2(_13681_),
    .B1_N(_13677_),
    .X(_13908_));
 sky130_fd_sc_hd__xnor2_1 _20632_ (.A(_13907_),
    .B(_13908_),
    .Y(_13909_));
 sky130_fd_sc_hd__and2_1 _20633_ (.A(_13896_),
    .B(_13909_),
    .X(_13910_));
 sky130_fd_sc_hd__nor2_1 _20634_ (.A(_13896_),
    .B(_13909_),
    .Y(_13911_));
 sky130_fd_sc_hd__or2_4 _20635_ (.A(_13910_),
    .B(_13911_),
    .X(_13912_));
 sky130_fd_sc_hd__nand2_2 _20636_ (.A(_13692_),
    .B(_13694_),
    .Y(_13913_));
 sky130_fd_sc_hd__o21ba_1 _20637_ (.A1(_13712_),
    .A2(_13717_),
    .B1_N(_13714_),
    .X(_13914_));
 sky130_fd_sc_hd__a22oi_1 _20638_ (.A1(_11664_),
    .A2(_13690_),
    .B1(_11666_),
    .B2(_11491_),
    .Y(_13915_));
 sky130_fd_sc_hd__and4_1 _20639_ (.A(_11825_),
    .B(_11656_),
    .C(_11599_),
    .D(_11927_),
    .X(_13916_));
 sky130_fd_sc_hd__nor2_2 _20640_ (.A(_13915_),
    .B(_13916_),
    .Y(_13917_));
 sky130_fd_sc_hd__clkbuf_2 _20641_ (.A(_12285_),
    .X(_13918_));
 sky130_fd_sc_hd__clkbuf_4 _20642_ (.A(_13918_),
    .X(_13919_));
 sky130_fd_sc_hd__nand2_2 _20643_ (.A(_11445_),
    .B(_13919_),
    .Y(_13920_));
 sky130_fd_sc_hd__xnor2_4 _20644_ (.A(_13917_),
    .B(_13920_),
    .Y(_13921_));
 sky130_fd_sc_hd__xnor2_1 _20645_ (.A(_13914_),
    .B(_13921_),
    .Y(_13922_));
 sky130_fd_sc_hd__xnor2_1 _20646_ (.A(_13913_),
    .B(_13922_),
    .Y(_13923_));
 sky130_fd_sc_hd__a21oi_1 _20647_ (.A1(_13697_),
    .A2(_13699_),
    .B1(_13923_),
    .Y(_13924_));
 sky130_fd_sc_hd__and3_1 _20648_ (.A(_13697_),
    .B(_13699_),
    .C(_13923_),
    .X(_13925_));
 sky130_fd_sc_hd__nor3_1 _20649_ (.A(_13912_),
    .B(_13924_),
    .C(_13925_),
    .Y(_13926_));
 sky130_fd_sc_hd__o21a_1 _20650_ (.A1(_13924_),
    .A2(_13925_),
    .B1(_13912_),
    .X(_13927_));
 sky130_fd_sc_hd__a211oi_1 _20651_ (.A1(_13886_),
    .A2(_13734_),
    .B1(_13926_),
    .C1(_13927_),
    .Y(_13928_));
 sky130_fd_sc_hd__o211a_1 _20652_ (.A1(_13926_),
    .A2(_13927_),
    .B1(_13886_),
    .C1(_13734_),
    .X(_13929_));
 sky130_fd_sc_hd__nor2_1 _20653_ (.A(_13928_),
    .B(_13929_),
    .Y(_13930_));
 sky130_fd_sc_hd__xnor2_2 _20654_ (.A(_13885_),
    .B(_13930_),
    .Y(_13931_));
 sky130_fd_sc_hd__nand2_1 _20655_ (.A(_13728_),
    .B(_13730_),
    .Y(_13932_));
 sky130_fd_sc_hd__nand2_1 _20656_ (.A(_11382_),
    .B(_11771_),
    .Y(_13933_));
 sky130_fd_sc_hd__clkbuf_2 _20657_ (.A(_12021_),
    .X(_13934_));
 sky130_fd_sc_hd__and4_1 _20658_ (.A(_11172_),
    .B(_11373_),
    .C(_11896_),
    .D(_13934_),
    .X(_13935_));
 sky130_fd_sc_hd__clkbuf_4 _20659_ (.A(_13713_),
    .X(_13936_));
 sky130_fd_sc_hd__clkbuf_4 _20660_ (.A(_12021_),
    .X(_13937_));
 sky130_fd_sc_hd__a22oi_1 _20661_ (.A1(_11278_),
    .A2(_13936_),
    .B1(_13937_),
    .B2(_11262_),
    .Y(_13938_));
 sky130_fd_sc_hd__nor2_1 _20662_ (.A(_13935_),
    .B(_13938_),
    .Y(_13939_));
 sky130_fd_sc_hd__xnor2_2 _20663_ (.A(_13933_),
    .B(_13939_),
    .Y(_13940_));
 sky130_fd_sc_hd__nand2_1 _20664_ (.A(_11161_),
    .B(_13720_),
    .Y(_13941_));
 sky130_fd_sc_hd__clkbuf_4 _20665_ (.A(_12328_),
    .X(_13942_));
 sky130_fd_sc_hd__and4_1 _20666_ (.A(_11037_),
    .B(_11039_),
    .C(_13942_),
    .D(_13721_),
    .X(_13943_));
 sky130_fd_sc_hd__clkbuf_2 _20667_ (.A(_12600_),
    .X(_13944_));
 sky130_fd_sc_hd__buf_4 _20668_ (.A(_13944_),
    .X(_13945_));
 sky130_fd_sc_hd__a22oi_2 _20669_ (.A1(_11270_),
    .A2(_12324_),
    .B1(_13945_),
    .B2(_11167_),
    .Y(_13946_));
 sky130_fd_sc_hd__nor2_1 _20670_ (.A(_13943_),
    .B(_13946_),
    .Y(_13947_));
 sky130_fd_sc_hd__xnor2_2 _20671_ (.A(_13941_),
    .B(_13947_),
    .Y(_13948_));
 sky130_fd_sc_hd__and2_1 _20672_ (.A(_13722_),
    .B(_13725_),
    .X(_13949_));
 sky130_fd_sc_hd__xnor2_1 _20673_ (.A(_13948_),
    .B(_13949_),
    .Y(_13950_));
 sky130_fd_sc_hd__xnor2_1 _20674_ (.A(_13940_),
    .B(_13950_),
    .Y(_13951_));
 sky130_fd_sc_hd__a21oi_1 _20675_ (.A1(_13748_),
    .A2(_13750_),
    .B1(_13951_),
    .Y(_13952_));
 sky130_fd_sc_hd__nand3_1 _20676_ (.A(_13748_),
    .B(_13750_),
    .C(_13951_),
    .Y(_13953_));
 sky130_fd_sc_hd__or2b_1 _20677_ (.A(_13952_),
    .B_N(_13953_),
    .X(_13954_));
 sky130_fd_sc_hd__xnor2_2 _20678_ (.A(_13932_),
    .B(_13954_),
    .Y(_13955_));
 sky130_fd_sc_hd__nand2_1 _20679_ (.A(_13742_),
    .B(_13746_),
    .Y(_13956_));
 sky130_fd_sc_hd__and2_1 _20680_ (.A(_13763_),
    .B(_13767_),
    .X(_13957_));
 sky130_fd_sc_hd__and4_1 _20681_ (.A(_11193_),
    .B(_11405_),
    .C(_13739_),
    .D(_13741_),
    .X(_13958_));
 sky130_fd_sc_hd__buf_2 _20682_ (.A(_11059_),
    .X(_13959_));
 sky130_fd_sc_hd__buf_2 _20683_ (.A(_13061_),
    .X(_13960_));
 sky130_fd_sc_hd__clkbuf_4 _20684_ (.A(_13960_),
    .X(_13961_));
 sky130_fd_sc_hd__a22oi_2 _20685_ (.A1(_13959_),
    .A2(_12772_),
    .B1(_13961_),
    .B2(_12361_),
    .Y(_13962_));
 sky130_fd_sc_hd__and4bb_1 _20686_ (.A_N(_13958_),
    .B_N(_13962_),
    .C(_11050_),
    .D(_12586_),
    .X(_13963_));
 sky130_fd_sc_hd__o2bb2a_1 _20687_ (.A1_N(_11050_),
    .A2_N(_12586_),
    .B1(_13958_),
    .B2(_13962_),
    .X(_13964_));
 sky130_fd_sc_hd__nor2_1 _20688_ (.A(_13963_),
    .B(_13964_),
    .Y(_13965_));
 sky130_fd_sc_hd__xnor2_2 _20689_ (.A(_13957_),
    .B(_13965_),
    .Y(_13966_));
 sky130_fd_sc_hd__xor2_2 _20690_ (.A(_13956_),
    .B(_13966_),
    .X(_13967_));
 sky130_fd_sc_hd__nand2_1 _20691_ (.A(_11343_),
    .B(_13055_),
    .Y(_13968_));
 sky130_fd_sc_hd__and4_1 _20692_ (.A(_10650_),
    .B(_10797_),
    .C(_13764_),
    .D(_13765_),
    .X(_13969_));
 sky130_fd_sc_hd__clkbuf_4 _20693_ (.A(_13760_),
    .X(_13970_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20694_ (.A(\genblk1.pcpi_mul.rs2[29] ),
    .X(_13971_));
 sky130_fd_sc_hd__clkbuf_4 _20695_ (.A(_13971_),
    .X(_13972_));
 sky130_fd_sc_hd__a22oi_2 _20696_ (.A1(_10666_),
    .A2(_13970_),
    .B1(_13972_),
    .B2(_10676_),
    .Y(_13973_));
 sky130_fd_sc_hd__nor2_1 _20697_ (.A(_13969_),
    .B(_13973_),
    .Y(_13974_));
 sky130_fd_sc_hd__xnor2_2 _20698_ (.A(_13968_),
    .B(_13974_),
    .Y(_13975_));
 sky130_fd_sc_hd__nand2_1 _20699_ (.A(_10630_),
    .B(_13752_),
    .Y(_13976_));
 sky130_fd_sc_hd__nand2_1 _20700_ (.A(_10635_),
    .B(_13756_),
    .Y(_13977_));
 sky130_fd_sc_hd__and2b_1 _20701_ (.A_N(_10710_),
    .B(_13802_),
    .X(_13978_));
 sky130_fd_sc_hd__xnor2_2 _20702_ (.A(_13977_),
    .B(_13978_),
    .Y(_13979_));
 sky130_fd_sc_hd__xnor2_2 _20703_ (.A(_13976_),
    .B(_13979_),
    .Y(_13980_));
 sky130_fd_sc_hd__xor2_2 _20704_ (.A(_13758_),
    .B(_13980_),
    .X(_13981_));
 sky130_fd_sc_hd__xnor2_2 _20705_ (.A(_13975_),
    .B(_13981_),
    .Y(_13982_));
 sky130_fd_sc_hd__xor2_2 _20706_ (.A(_13769_),
    .B(_13982_),
    .X(_13983_));
 sky130_fd_sc_hd__xnor2_2 _20707_ (.A(_13967_),
    .B(_13983_),
    .Y(_13984_));
 sky130_fd_sc_hd__nand2_1 _20708_ (.A(_13771_),
    .B(_13773_),
    .Y(_13985_));
 sky130_fd_sc_hd__xnor2_2 _20709_ (.A(_13984_),
    .B(_13985_),
    .Y(_13986_));
 sky130_fd_sc_hd__xnor2_2 _20710_ (.A(_13955_),
    .B(_13986_),
    .Y(_13987_));
 sky130_fd_sc_hd__nand2_1 _20711_ (.A(_13775_),
    .B(_13777_),
    .Y(_13988_));
 sky130_fd_sc_hd__xnor2_2 _20712_ (.A(_13987_),
    .B(_13988_),
    .Y(_13989_));
 sky130_fd_sc_hd__xor2_2 _20713_ (.A(_13931_),
    .B(_13989_),
    .X(_13990_));
 sky130_fd_sc_hd__or2_1 _20714_ (.A(_13779_),
    .B(_13781_),
    .X(_13991_));
 sky130_fd_sc_hd__xor2_2 _20715_ (.A(_13990_),
    .B(_13991_),
    .X(_13992_));
 sky130_fd_sc_hd__xnor2_1 _20716_ (.A(_13884_),
    .B(_13992_),
    .Y(_13993_));
 sky130_fd_sc_hd__nand2_1 _20717_ (.A(_13783_),
    .B(_13785_),
    .Y(_13994_));
 sky130_fd_sc_hd__xnor2_1 _20718_ (.A(_13993_),
    .B(_13994_),
    .Y(_13995_));
 sky130_fd_sc_hd__xnor2_1 _20719_ (.A(_13810_),
    .B(_13995_),
    .Y(_13996_));
 sky130_fd_sc_hd__nor2_1 _20720_ (.A(_13787_),
    .B(_13789_),
    .Y(_13997_));
 sky130_fd_sc_hd__xnor2_2 _20721_ (.A(_13996_),
    .B(_13997_),
    .Y(_13998_));
 sky130_fd_sc_hd__xnor2_4 _20722_ (.A(_13801_),
    .B(_13998_),
    .Y(_13999_));
 sky130_fd_sc_hd__nor2_2 _20723_ (.A(_13791_),
    .B(_13793_),
    .Y(_14000_));
 sky130_fd_sc_hd__xor2_4 _20724_ (.A(_13999_),
    .B(_14000_),
    .X(_14001_));
 sky130_fd_sc_hd__or2_1 _20725_ (.A(_13799_),
    .B(_13796_),
    .X(_14002_));
 sky130_fd_sc_hd__and4bb_1 _20726_ (.A_N(_13261_),
    .B_N(_13429_),
    .C(_13590_),
    .D(_13798_),
    .X(_14003_));
 sky130_fd_sc_hd__o31ai_1 _20727_ (.A1(_12812_),
    .A2(_12957_),
    .A3(_13262_),
    .B1(_13264_),
    .Y(_14004_));
 sky130_fd_sc_hd__nand2_1 _20728_ (.A(_13590_),
    .B(_13798_),
    .Y(_14005_));
 sky130_fd_sc_hd__o2bb2a_2 _20729_ (.A1_N(_14003_),
    .A2_N(_14004_),
    .B1(_13592_),
    .B2(_14005_),
    .X(_14006_));
 sky130_fd_sc_hd__and3_4 _20730_ (.A(_13797_),
    .B(_14002_),
    .C(_14006_),
    .X(_14007_));
 sky130_fd_sc_hd__or4b_4 _20731_ (.A(_12666_),
    .B(_12956_),
    .C(_13262_),
    .D_N(_14003_),
    .X(_14008_));
 sky130_fd_sc_hd__a21o_4 _20732_ (.A1(_12668_),
    .A2(_12673_),
    .B1(_14008_),
    .X(_14009_));
 sky130_fd_sc_hd__nand2_2 _20733_ (.A(_14007_),
    .B(_14009_),
    .Y(_14010_));
 sky130_fd_sc_hd__xor2_4 _20734_ (.A(_14001_),
    .B(_14010_),
    .X(_00078_));
 sky130_fd_sc_hd__nor2_1 _20735_ (.A(_13999_),
    .B(_14000_),
    .Y(_14011_));
 sky130_fd_sc_hd__a21oi_2 _20736_ (.A1(_14001_),
    .A2(_14010_),
    .B1(_14011_),
    .Y(_14012_));
 sky130_fd_sc_hd__or2b_1 _20737_ (.A(_13997_),
    .B_N(_13996_),
    .X(_14013_));
 sky130_fd_sc_hd__nand2_1 _20738_ (.A(_13801_),
    .B(_13998_),
    .Y(_14014_));
 sky130_fd_sc_hd__a21o_1 _20739_ (.A1(_13805_),
    .A2(_13809_),
    .B1(_13807_),
    .X(_14015_));
 sky130_fd_sc_hd__and2b_1 _20740_ (.A_N(_13883_),
    .B(_13811_),
    .X(_14016_));
 sky130_fd_sc_hd__a21o_1 _20741_ (.A1(_13812_),
    .A2(_13882_),
    .B1(_14016_),
    .X(_14017_));
 sky130_fd_sc_hd__nor2_1 _20742_ (.A(_13850_),
    .B(_13852_),
    .Y(_14018_));
 sky130_fd_sc_hd__xnor2_2 _20743_ (.A(_14017_),
    .B(_14018_),
    .Y(_14019_));
 sky130_fd_sc_hd__or2_2 _20744_ (.A(_13878_),
    .B(_13880_),
    .X(_14020_));
 sky130_fd_sc_hd__o21ba_1 _20745_ (.A1(_13885_),
    .A2(_13929_),
    .B1_N(_13928_),
    .X(_14021_));
 sky130_fd_sc_hd__and2b_1 _20746_ (.A_N(_13845_),
    .B(_13844_),
    .X(_14022_));
 sky130_fd_sc_hd__buf_2 _20747_ (.A(_13817_),
    .X(_14023_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20748_ (.A(\genblk1.pcpi_mul.rs1[32] ),
    .X(_14024_));
 sky130_fd_sc_hd__and3_2 _20749_ (.A(_11044_),
    .B(_11041_),
    .C(_14024_),
    .X(_14025_));
 sky130_fd_sc_hd__buf_2 _20750_ (.A(_14024_),
    .X(_14026_));
 sky130_fd_sc_hd__a22oi_1 _20751_ (.A1(_10612_),
    .A2(_13830_),
    .B1(_14026_),
    .B2(_10627_),
    .Y(_14027_));
 sky130_fd_sc_hd__a21oi_1 _20752_ (.A1(_13831_),
    .A2(_14025_),
    .B1(_14027_),
    .Y(_14028_));
 sky130_fd_sc_hd__a21oi_1 _20753_ (.A1(_11368_),
    .A2(_14023_),
    .B1(_14028_),
    .Y(_14029_));
 sky130_fd_sc_hd__and3_1 _20754_ (.A(_10680_),
    .B(_13817_),
    .C(_14028_),
    .X(_14030_));
 sky130_fd_sc_hd__or2_1 _20755_ (.A(_14029_),
    .B(_14030_),
    .X(_14031_));
 sky130_fd_sc_hd__a22oi_1 _20756_ (.A1(_11385_),
    .A2(_13836_),
    .B1(_13814_),
    .B2(_11387_),
    .Y(_14032_));
 sky130_fd_sc_hd__clkbuf_2 _20757_ (.A(_13292_),
    .X(_14033_));
 sky130_fd_sc_hd__and4_1 _20758_ (.A(_10672_),
    .B(_11282_),
    .C(_13839_),
    .D(_14033_),
    .X(_14034_));
 sky130_fd_sc_hd__nor2_1 _20759_ (.A(_14032_),
    .B(_14034_),
    .Y(_14035_));
 sky130_fd_sc_hd__xnor2_1 _20760_ (.A(_13843_),
    .B(_14035_),
    .Y(_14036_));
 sky130_fd_sc_hd__buf_2 _20761_ (.A(_14024_),
    .X(_14037_));
 sky130_fd_sc_hd__buf_2 _20762_ (.A(_14037_),
    .X(_14038_));
 sky130_fd_sc_hd__a31o_1 _20763_ (.A1(_10584_),
    .A2(_14038_),
    .A3(_13841_),
    .B1(_13840_),
    .X(_14039_));
 sky130_fd_sc_hd__xnor2_1 _20764_ (.A(_14036_),
    .B(_14039_),
    .Y(_14040_));
 sky130_fd_sc_hd__xor2_1 _20765_ (.A(_14031_),
    .B(_14040_),
    .X(_14041_));
 sky130_fd_sc_hd__o21a_4 _20766_ (.A1(_14022_),
    .A2(_13847_),
    .B1(_14041_),
    .X(_14042_));
 sky130_fd_sc_hd__nor3_1 _20767_ (.A(_14022_),
    .B(_13847_),
    .C(_14041_),
    .Y(_14043_));
 sky130_fd_sc_hd__or2_1 _20768_ (.A(_14042_),
    .B(_14043_),
    .X(_14044_));
 sky130_fd_sc_hd__a21oi_4 _20769_ (.A1(_13832_),
    .A2(_13834_),
    .B1(_14044_),
    .Y(_14045_));
 sky130_fd_sc_hd__and3_2 _20770_ (.A(_13832_),
    .B(_13834_),
    .C(_14044_),
    .X(_14046_));
 sky130_fd_sc_hd__nor2_1 _20771_ (.A(_14045_),
    .B(_14046_),
    .Y(_14047_));
 sky130_vsdinv _20772_ (.A(_13874_),
    .Y(_14048_));
 sky130_fd_sc_hd__or2b_1 _20773_ (.A(_13857_),
    .B_N(_13871_),
    .X(_14049_));
 sky130_fd_sc_hd__nand2_4 _20774_ (.A(_13856_),
    .B(_13872_),
    .Y(_14050_));
 sky130_fd_sc_hd__and2b_1 _20775_ (.A_N(_13908_),
    .B(_13907_),
    .X(_14051_));
 sky130_fd_sc_hd__o21ba_1 _20776_ (.A1(_13862_),
    .A2(_13870_),
    .B1_N(_13865_),
    .X(_14052_));
 sky130_fd_sc_hd__o21ba_1 _20777_ (.A1(_13889_),
    .A2(_13894_),
    .B1_N(_13892_),
    .X(_14053_));
 sky130_fd_sc_hd__a22oi_1 _20778_ (.A1(_13858_),
    .A2(_13864_),
    .B1(_13286_),
    .B2(_10784_),
    .Y(_14054_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20779_ (.A(_11086_),
    .X(_14055_));
 sky130_fd_sc_hd__clkbuf_2 _20780_ (.A(_12973_),
    .X(_14056_));
 sky130_fd_sc_hd__and4_1 _20781_ (.A(_13863_),
    .B(_14055_),
    .C(_13637_),
    .D(_14056_),
    .X(_14057_));
 sky130_fd_sc_hd__nor2_1 _20782_ (.A(_14054_),
    .B(_14057_),
    .Y(_14058_));
 sky130_fd_sc_hd__buf_2 _20783_ (.A(_13446_),
    .X(_14059_));
 sky130_fd_sc_hd__nand2_1 _20784_ (.A(_11080_),
    .B(_14059_),
    .Y(_14060_));
 sky130_fd_sc_hd__xnor2_1 _20785_ (.A(_14058_),
    .B(_14060_),
    .Y(_14061_));
 sky130_fd_sc_hd__xnor2_1 _20786_ (.A(_14053_),
    .B(_14061_),
    .Y(_14062_));
 sky130_fd_sc_hd__xnor2_1 _20787_ (.A(_14052_),
    .B(_14062_),
    .Y(_14063_));
 sky130_fd_sc_hd__o21a_1 _20788_ (.A1(_14051_),
    .A2(_13910_),
    .B1(_14063_),
    .X(_14064_));
 sky130_fd_sc_hd__nor3_1 _20789_ (.A(_14051_),
    .B(_13910_),
    .C(_14063_),
    .Y(_14065_));
 sky130_fd_sc_hd__a211oi_4 _20790_ (.A1(_14049_),
    .A2(_14050_),
    .B1(_14064_),
    .C1(net360),
    .Y(_14066_));
 sky130_fd_sc_hd__o211a_2 _20791_ (.A1(_14064_),
    .A2(_14065_),
    .B1(_14049_),
    .C1(_14050_),
    .X(_14067_));
 sky130_fd_sc_hd__a211o_1 _20792_ (.A1(_14048_),
    .A2(_13876_),
    .B1(_14066_),
    .C1(_14067_),
    .X(_14068_));
 sky130_fd_sc_hd__o211ai_1 _20793_ (.A1(_14066_),
    .A2(_14067_),
    .B1(_14048_),
    .C1(_13876_),
    .Y(_14069_));
 sky130_fd_sc_hd__nand2_1 _20794_ (.A(_14068_),
    .B(_14069_),
    .Y(_14070_));
 sky130_fd_sc_hd__xnor2_2 _20795_ (.A(_14047_),
    .B(_14070_),
    .Y(_14071_));
 sky130_fd_sc_hd__xnor2_2 _20796_ (.A(_14021_),
    .B(_14071_),
    .Y(_14072_));
 sky130_fd_sc_hd__xor2_2 _20797_ (.A(_14020_),
    .B(_14072_),
    .X(_14073_));
 sky130_fd_sc_hd__or2_1 _20798_ (.A(_13924_),
    .B(_13926_),
    .X(_14074_));
 sky130_fd_sc_hd__a21o_1 _20799_ (.A1(_13932_),
    .A2(_13953_),
    .B1(_13952_),
    .X(_14075_));
 sky130_fd_sc_hd__buf_2 _20800_ (.A(_12690_),
    .X(_14076_));
 sky130_fd_sc_hd__buf_2 _20801_ (.A(_14076_),
    .X(_14077_));
 sky130_fd_sc_hd__nand2_1 _20802_ (.A(_11138_),
    .B(_14077_),
    .Y(_14078_));
 sky130_fd_sc_hd__and4_1 _20803_ (.A(_13669_),
    .B(_11112_),
    .C(_12694_),
    .D(_13887_),
    .X(_14079_));
 sky130_fd_sc_hd__buf_2 _20804_ (.A(_12538_),
    .X(_14080_));
 sky130_fd_sc_hd__buf_2 _20805_ (.A(_14080_),
    .X(_14081_));
 sky130_fd_sc_hd__a22oi_1 _20806_ (.A1(_13665_),
    .A2(_13891_),
    .B1(_14081_),
    .B2(_13670_),
    .Y(_14082_));
 sky130_fd_sc_hd__nor2_1 _20807_ (.A(_14079_),
    .B(_14082_),
    .Y(_14083_));
 sky130_fd_sc_hd__xnor2_1 _20808_ (.A(_14078_),
    .B(_14083_),
    .Y(_14084_));
 sky130_fd_sc_hd__nand2_1 _20809_ (.A(_11136_),
    .B(_13668_),
    .Y(_14085_));
 sky130_fd_sc_hd__clkbuf_2 _20810_ (.A(_11356_),
    .X(_14086_));
 sky130_fd_sc_hd__buf_2 _20811_ (.A(_11458_),
    .X(_14087_));
 sky130_fd_sc_hd__and4_1 _20812_ (.A(_14086_),
    .B(_14087_),
    .C(_11959_),
    .D(_12145_),
    .X(_14088_));
 sky130_fd_sc_hd__a22oi_2 _20813_ (.A1(_13903_),
    .A2(_13901_),
    .B1(_13663_),
    .B2(_13899_),
    .Y(_14089_));
 sky130_fd_sc_hd__nor2_1 _20814_ (.A(_14088_),
    .B(_14089_),
    .Y(_14090_));
 sky130_fd_sc_hd__xnor2_1 _20815_ (.A(_14085_),
    .B(_14090_),
    .Y(_14091_));
 sky130_fd_sc_hd__o21ba_1 _20816_ (.A1(_13898_),
    .A2(_13905_),
    .B1_N(_13902_),
    .X(_14092_));
 sky130_fd_sc_hd__xnor2_1 _20817_ (.A(_14091_),
    .B(_14092_),
    .Y(_14093_));
 sky130_fd_sc_hd__and2_1 _20818_ (.A(_14084_),
    .B(_14093_),
    .X(_14094_));
 sky130_fd_sc_hd__nor2_1 _20819_ (.A(_14084_),
    .B(_14093_),
    .Y(_14095_));
 sky130_fd_sc_hd__or2_2 _20820_ (.A(_14094_),
    .B(_14095_),
    .X(_14096_));
 sky130_fd_sc_hd__or2b_1 _20821_ (.A(_13914_),
    .B_N(_13921_),
    .X(_14097_));
 sky130_fd_sc_hd__nand2_1 _20822_ (.A(_13913_),
    .B(_13922_),
    .Y(_14098_));
 sky130_fd_sc_hd__buf_2 _20823_ (.A(_11561_),
    .X(_14099_));
 sky130_fd_sc_hd__a31o_2 _20824_ (.A1(_14099_),
    .A2(_13919_),
    .A3(_13917_),
    .B1(_13916_),
    .X(_14100_));
 sky130_fd_sc_hd__o21ba_1 _20825_ (.A1(_13933_),
    .A2(_13938_),
    .B1_N(_13935_),
    .X(_14101_));
 sky130_fd_sc_hd__nand2_1 _20826_ (.A(_11775_),
    .B(_13904_),
    .Y(_14102_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20827_ (.A(_11662_),
    .X(_14103_));
 sky130_fd_sc_hd__and4_1 _20828_ (.A(_14103_),
    .B(_13689_),
    .C(_11665_),
    .D(_11708_),
    .X(_14104_));
 sky130_fd_sc_hd__buf_2 _20829_ (.A(_11923_),
    .X(_14105_));
 sky130_fd_sc_hd__a22oi_1 _20830_ (.A1(_13695_),
    .A2(_11927_),
    .B1(_11820_),
    .B2(_14105_),
    .Y(_14106_));
 sky130_fd_sc_hd__nor2_1 _20831_ (.A(_14104_),
    .B(_14106_),
    .Y(_14107_));
 sky130_fd_sc_hd__xnor2_2 _20832_ (.A(_14102_),
    .B(_14107_),
    .Y(_14108_));
 sky130_fd_sc_hd__xnor2_2 _20833_ (.A(_14101_),
    .B(_14108_),
    .Y(_14109_));
 sky130_fd_sc_hd__xnor2_2 _20834_ (.A(_14100_),
    .B(_14109_),
    .Y(_14110_));
 sky130_fd_sc_hd__a21oi_1 _20835_ (.A1(_14097_),
    .A2(_14098_),
    .B1(_14110_),
    .Y(_14111_));
 sky130_fd_sc_hd__and3_1 _20836_ (.A(_14097_),
    .B(_14098_),
    .C(_14110_),
    .X(_14112_));
 sky130_fd_sc_hd__nor3_1 _20837_ (.A(_14096_),
    .B(_14111_),
    .C(_14112_),
    .Y(_14113_));
 sky130_fd_sc_hd__o21a_1 _20838_ (.A1(_14111_),
    .A2(_14112_),
    .B1(_14096_),
    .X(_14114_));
 sky130_fd_sc_hd__or2_1 _20839_ (.A(_14113_),
    .B(_14114_),
    .X(_14115_));
 sky130_fd_sc_hd__xnor2_2 _20840_ (.A(_14075_),
    .B(_14115_),
    .Y(_14116_));
 sky130_fd_sc_hd__xor2_2 _20841_ (.A(_14074_),
    .B(_14116_),
    .X(_14117_));
 sky130_fd_sc_hd__and2b_1 _20842_ (.A_N(_13949_),
    .B(_13948_),
    .X(_14118_));
 sky130_fd_sc_hd__a21o_1 _20843_ (.A1(_13940_),
    .A2(_13950_),
    .B1(_14118_),
    .X(_14119_));
 sky130_fd_sc_hd__or3_1 _20844_ (.A(_13957_),
    .B(_13963_),
    .C(_13964_),
    .X(_14120_));
 sky130_fd_sc_hd__nand2_1 _20845_ (.A(_13956_),
    .B(_13966_),
    .Y(_14121_));
 sky130_fd_sc_hd__nand2_1 _20846_ (.A(_11826_),
    .B(_12591_),
    .Y(_14122_));
 sky130_fd_sc_hd__clkbuf_2 _20847_ (.A(_12235_),
    .X(_14123_));
 sky130_fd_sc_hd__and4_1 _20848_ (.A(_11479_),
    .B(_11482_),
    .C(_14123_),
    .D(_13934_),
    .X(_14124_));
 sky130_fd_sc_hd__a22oi_2 _20849_ (.A1(_11477_),
    .A2(_11891_),
    .B1(_13937_),
    .B2(_11278_),
    .Y(_14125_));
 sky130_fd_sc_hd__nor2_1 _20850_ (.A(_14124_),
    .B(_14125_),
    .Y(_14126_));
 sky130_fd_sc_hd__xnor2_1 _20851_ (.A(_14122_),
    .B(_14126_),
    .Y(_14127_));
 sky130_fd_sc_hd__nand2_1 _20852_ (.A(_11474_),
    .B(_13720_),
    .Y(_14128_));
 sky130_fd_sc_hd__buf_2 _20853_ (.A(_13376_),
    .X(_14129_));
 sky130_fd_sc_hd__and4_1 _20854_ (.A(_11156_),
    .B(_11264_),
    .C(_12329_),
    .D(_14129_),
    .X(_14130_));
 sky130_fd_sc_hd__clkbuf_2 _20855_ (.A(_12327_),
    .X(_14131_));
 sky130_fd_sc_hd__clkbuf_4 _20856_ (.A(_14131_),
    .X(_14132_));
 sky130_fd_sc_hd__a22oi_4 _20857_ (.A1(_11068_),
    .A2(_14132_),
    .B1(_13945_),
    .B2(_11039_),
    .Y(_14133_));
 sky130_fd_sc_hd__nor2_1 _20858_ (.A(_14130_),
    .B(_14133_),
    .Y(_14134_));
 sky130_fd_sc_hd__xnor2_1 _20859_ (.A(_14128_),
    .B(_14134_),
    .Y(_14135_));
 sky130_fd_sc_hd__o21ba_1 _20860_ (.A1(_13941_),
    .A2(_13946_),
    .B1_N(_13943_),
    .X(_14136_));
 sky130_fd_sc_hd__xnor2_1 _20861_ (.A(_14135_),
    .B(_14136_),
    .Y(_14137_));
 sky130_fd_sc_hd__xnor2_1 _20862_ (.A(_14127_),
    .B(_14137_),
    .Y(_14138_));
 sky130_fd_sc_hd__a21oi_1 _20863_ (.A1(_14120_),
    .A2(_14121_),
    .B1(_14138_),
    .Y(_14139_));
 sky130_fd_sc_hd__and3_1 _20864_ (.A(_14120_),
    .B(_14121_),
    .C(_14138_),
    .X(_14140_));
 sky130_fd_sc_hd__nor2_1 _20865_ (.A(_14139_),
    .B(_14140_),
    .Y(_14141_));
 sky130_fd_sc_hd__xor2_2 _20866_ (.A(_14119_),
    .B(_14141_),
    .X(_14142_));
 sky130_fd_sc_hd__o21ba_1 _20867_ (.A1(_13968_),
    .A2(_13973_),
    .B1_N(_13969_),
    .X(_14143_));
 sky130_fd_sc_hd__and4_2 _20868_ (.A(_11062_),
    .B(_11175_),
    .C(_13558_),
    .D(_13556_),
    .X(_14144_));
 sky130_fd_sc_hd__a22oi_2 _20869_ (.A1(_11177_),
    .A2(_12771_),
    .B1(_13960_),
    .B2(_10973_),
    .Y(_14145_));
 sky130_fd_sc_hd__and4bb_1 _20870_ (.A_N(_14144_),
    .B_N(_14145_),
    .C(_11386_),
    .D(_12585_),
    .X(_14146_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20871_ (.A(_12584_),
    .X(_14147_));
 sky130_fd_sc_hd__o2bb2a_1 _20872_ (.A1_N(_11386_),
    .A2_N(_14147_),
    .B1(_14144_),
    .B2(_14145_),
    .X(_14148_));
 sky130_fd_sc_hd__nor2_1 _20873_ (.A(_14146_),
    .B(_14148_),
    .Y(_14149_));
 sky130_fd_sc_hd__xnor2_1 _20874_ (.A(_14143_),
    .B(_14149_),
    .Y(_14150_));
 sky130_fd_sc_hd__o21ai_1 _20875_ (.A1(_13958_),
    .A2(_13963_),
    .B1(_14150_),
    .Y(_14151_));
 sky130_fd_sc_hd__or3_1 _20876_ (.A(_13958_),
    .B(_13963_),
    .C(_14150_),
    .X(_14152_));
 sky130_fd_sc_hd__and2_1 _20877_ (.A(_14151_),
    .B(_14152_),
    .X(_14153_));
 sky130_fd_sc_hd__clkbuf_2 _20878_ (.A(_13054_),
    .X(_14154_));
 sky130_fd_sc_hd__nand2_1 _20879_ (.A(_11404_),
    .B(_14154_),
    .Y(_14155_));
 sky130_fd_sc_hd__and4_1 _20880_ (.A(_10797_),
    .B(_11199_),
    .C(_13223_),
    .D(_13971_),
    .X(_14156_));
 sky130_fd_sc_hd__a22oi_2 _20881_ (.A1(_11091_),
    .A2(_13761_),
    .B1(_13762_),
    .B2(_10666_),
    .Y(_14157_));
 sky130_fd_sc_hd__nor2_1 _20882_ (.A(_14156_),
    .B(_14157_),
    .Y(_14158_));
 sky130_fd_sc_hd__xnor2_2 _20883_ (.A(_14155_),
    .B(_14158_),
    .Y(_14159_));
 sky130_fd_sc_hd__buf_2 _20884_ (.A(\genblk1.pcpi_mul.rs2[30] ),
    .X(_14160_));
 sky130_fd_sc_hd__nand2_1 _20885_ (.A(_10676_),
    .B(_14160_),
    .Y(_14161_));
 sky130_fd_sc_hd__and2b_1 _20886_ (.A_N(_10594_),
    .B(_13802_),
    .X(_14162_));
 sky130_fd_sc_hd__nand2_1 _20887_ (.A(_11777_),
    .B(_13756_),
    .Y(_14163_));
 sky130_fd_sc_hd__xnor2_2 _20888_ (.A(_14162_),
    .B(_14163_),
    .Y(_14164_));
 sky130_fd_sc_hd__xnor2_2 _20889_ (.A(_14161_),
    .B(_14164_),
    .Y(_14165_));
 sky130_fd_sc_hd__clkbuf_4 _20890_ (.A(_13541_),
    .X(_14166_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20891_ (.A(\genblk1.pcpi_mul.rs2[31] ),
    .X(_14167_));
 sky130_fd_sc_hd__buf_2 _20892_ (.A(_14167_),
    .X(_14168_));
 sky130_fd_sc_hd__and3_1 _20893_ (.A(_10638_),
    .B(_14168_),
    .C(_13978_),
    .X(_14169_));
 sky130_fd_sc_hd__a31o_1 _20894_ (.A1(_10609_),
    .A2(_14166_),
    .A3(_13979_),
    .B1(_14169_),
    .X(_14170_));
 sky130_fd_sc_hd__xor2_2 _20895_ (.A(_14165_),
    .B(_14170_),
    .X(_14171_));
 sky130_fd_sc_hd__xnor2_2 _20896_ (.A(_14159_),
    .B(_14171_),
    .Y(_14172_));
 sky130_fd_sc_hd__nand2_1 _20897_ (.A(_13758_),
    .B(_13980_),
    .Y(_14173_));
 sky130_fd_sc_hd__a21boi_2 _20898_ (.A1(_13975_),
    .A2(_13981_),
    .B1_N(_14173_),
    .Y(_14174_));
 sky130_fd_sc_hd__xnor2_1 _20899_ (.A(_14172_),
    .B(_14174_),
    .Y(_14175_));
 sky130_fd_sc_hd__xnor2_2 _20900_ (.A(_14153_),
    .B(_14175_),
    .Y(_14176_));
 sky130_fd_sc_hd__nor2_1 _20901_ (.A(_13769_),
    .B(_13982_),
    .Y(_14177_));
 sky130_fd_sc_hd__a21oi_2 _20902_ (.A1(_13967_),
    .A2(_13983_),
    .B1(_14177_),
    .Y(_14178_));
 sky130_fd_sc_hd__xnor2_2 _20903_ (.A(_14176_),
    .B(_14178_),
    .Y(_14179_));
 sky130_fd_sc_hd__xnor2_2 _20904_ (.A(_14142_),
    .B(_14179_),
    .Y(_14180_));
 sky130_fd_sc_hd__and2b_1 _20905_ (.A_N(_13984_),
    .B(_13985_),
    .X(_14181_));
 sky130_fd_sc_hd__a21oi_2 _20906_ (.A1(_13955_),
    .A2(_13986_),
    .B1(_14181_),
    .Y(_14182_));
 sky130_fd_sc_hd__xor2_2 _20907_ (.A(_14180_),
    .B(_14182_),
    .X(_14183_));
 sky130_fd_sc_hd__xnor2_2 _20908_ (.A(_14117_),
    .B(_14183_),
    .Y(_14184_));
 sky130_fd_sc_hd__and2b_1 _20909_ (.A_N(_13987_),
    .B(_13988_),
    .X(_14185_));
 sky130_fd_sc_hd__a21oi_2 _20910_ (.A1(_13931_),
    .A2(_13989_),
    .B1(_14185_),
    .Y(_14186_));
 sky130_fd_sc_hd__xor2_2 _20911_ (.A(_14184_),
    .B(_14186_),
    .X(_14187_));
 sky130_fd_sc_hd__xnor2_2 _20912_ (.A(_14073_),
    .B(_14187_),
    .Y(_14188_));
 sky130_fd_sc_hd__and2_1 _20913_ (.A(_13990_),
    .B(_13991_),
    .X(_14189_));
 sky130_fd_sc_hd__a21oi_2 _20914_ (.A1(_13884_),
    .A2(_13992_),
    .B1(_14189_),
    .Y(_14190_));
 sky130_fd_sc_hd__xor2_2 _20915_ (.A(_14188_),
    .B(_14190_),
    .X(_14191_));
 sky130_fd_sc_hd__xor2_2 _20916_ (.A(_14019_),
    .B(_14191_),
    .X(_14192_));
 sky130_vsdinv _20917_ (.A(_13810_),
    .Y(_14193_));
 sky130_fd_sc_hd__and2b_1 _20918_ (.A_N(_13993_),
    .B(_13994_),
    .X(_14194_));
 sky130_fd_sc_hd__a21oi_1 _20919_ (.A1(_14193_),
    .A2(_13995_),
    .B1(_14194_),
    .Y(_14195_));
 sky130_fd_sc_hd__xnor2_2 _20920_ (.A(_14192_),
    .B(_14195_),
    .Y(_14196_));
 sky130_fd_sc_hd__xnor2_1 _20921_ (.A(_14015_),
    .B(_14196_),
    .Y(_14197_));
 sky130_fd_sc_hd__nand3_1 _20922_ (.A(_14013_),
    .B(_14014_),
    .C(_14197_),
    .Y(_14198_));
 sky130_vsdinv _20923_ (.A(_14198_),
    .Y(_14199_));
 sky130_fd_sc_hd__a21oi_1 _20924_ (.A1(_14013_),
    .A2(_14014_),
    .B1(_14197_),
    .Y(_14200_));
 sky130_fd_sc_hd__nor2_2 _20925_ (.A(_14199_),
    .B(_14200_),
    .Y(_14201_));
 sky130_fd_sc_hd__xnor2_4 _20926_ (.A(_14012_),
    .B(_14201_),
    .Y(_00079_));
 sky130_fd_sc_hd__o21a_2 _20927_ (.A1(_13850_),
    .A2(_13852_),
    .B1(_14017_),
    .X(_14202_));
 sky130_fd_sc_hd__and2b_1 _20928_ (.A_N(_14021_),
    .B(_14071_),
    .X(_14203_));
 sky130_fd_sc_hd__a21o_2 _20929_ (.A1(_14020_),
    .A2(_14072_),
    .B1(_14203_),
    .X(_14204_));
 sky130_fd_sc_hd__nor2_2 _20930_ (.A(_14042_),
    .B(_14045_),
    .Y(_14205_));
 sky130_fd_sc_hd__xnor2_4 _20931_ (.A(_14204_),
    .B(_14205_),
    .Y(_14206_));
 sky130_fd_sc_hd__a21bo_2 _20932_ (.A1(_14047_),
    .A2(_14069_),
    .B1_N(_14068_),
    .X(_14207_));
 sky130_fd_sc_hd__or2b_1 _20933_ (.A(_14115_),
    .B_N(_14075_),
    .X(_14208_));
 sky130_fd_sc_hd__a21bo_1 _20934_ (.A1(_14074_),
    .A2(_14116_),
    .B1_N(_14208_),
    .X(_14209_));
 sky130_fd_sc_hd__buf_2 _20935_ (.A(_13618_),
    .X(_14210_));
 sky130_fd_sc_hd__clkbuf_2 _20936_ (.A(_14210_),
    .X(_14211_));
 sky130_fd_sc_hd__buf_2 _20937_ (.A(_14211_),
    .X(_14212_));
 sky130_fd_sc_hd__buf_2 _20938_ (.A(_14212_),
    .X(_14213_));
 sky130_fd_sc_hd__buf_2 _20939_ (.A(_14213_),
    .X(_14214_));
 sky130_fd_sc_hd__a21oi_4 _20940_ (.A1(_14214_),
    .A2(_14025_),
    .B1(_14030_),
    .Y(_14215_));
 sky130_fd_sc_hd__nand2_1 _20941_ (.A(_14036_),
    .B(_14039_),
    .Y(_14216_));
 sky130_fd_sc_hd__or2_2 _20942_ (.A(_14031_),
    .B(_14040_),
    .X(_14217_));
 sky130_fd_sc_hd__o21ai_1 _20943_ (.A1(_10641_),
    .A2(_10612_),
    .B1(_13842_),
    .Y(_14218_));
 sky130_fd_sc_hd__nor2_4 _20944_ (.A(_14025_),
    .B(_14218_),
    .Y(_14219_));
 sky130_fd_sc_hd__nand2_1 _20945_ (.A(_11368_),
    .B(_14212_),
    .Y(_14220_));
 sky130_fd_sc_hd__xor2_2 _20946_ (.A(_14219_),
    .B(_14220_),
    .X(_14221_));
 sky130_fd_sc_hd__buf_2 _20947_ (.A(_13843_),
    .X(_14222_));
 sky130_fd_sc_hd__buf_4 _20948_ (.A(_11282_),
    .X(_14223_));
 sky130_fd_sc_hd__a22oi_4 _20949_ (.A1(_14223_),
    .A2(_13814_),
    .B1(_13829_),
    .B2(_10663_),
    .Y(_14224_));
 sky130_fd_sc_hd__clkbuf_2 _20950_ (.A(_13605_),
    .X(_14225_));
 sky130_fd_sc_hd__and4_1 _20951_ (.A(_11387_),
    .B(_11385_),
    .C(_13824_),
    .D(_14225_),
    .X(_14226_));
 sky130_fd_sc_hd__nor2_1 _20952_ (.A(_14224_),
    .B(_14226_),
    .Y(_14227_));
 sky130_fd_sc_hd__xnor2_1 _20953_ (.A(_14222_),
    .B(_14227_),
    .Y(_14228_));
 sky130_fd_sc_hd__a31o_1 _20954_ (.A1(_10585_),
    .A2(_14038_),
    .A3(_14035_),
    .B1(_14034_),
    .X(_14229_));
 sky130_fd_sc_hd__xnor2_1 _20955_ (.A(_14228_),
    .B(_14229_),
    .Y(_14230_));
 sky130_fd_sc_hd__or2_1 _20956_ (.A(_14221_),
    .B(_14230_),
    .X(_14231_));
 sky130_fd_sc_hd__nand2_1 _20957_ (.A(_14221_),
    .B(_14230_),
    .Y(_14232_));
 sky130_fd_sc_hd__nand2_1 _20958_ (.A(_14231_),
    .B(_14232_),
    .Y(_14233_));
 sky130_fd_sc_hd__a21o_1 _20959_ (.A1(_14216_),
    .A2(_14217_),
    .B1(_14233_),
    .X(_14234_));
 sky130_fd_sc_hd__nand3_1 _20960_ (.A(_14216_),
    .B(_14217_),
    .C(_14233_),
    .Y(_14235_));
 sky130_fd_sc_hd__nand2_2 _20961_ (.A(_14234_),
    .B(_14235_),
    .Y(_14236_));
 sky130_fd_sc_hd__xor2_4 _20962_ (.A(_14215_),
    .B(_14236_),
    .X(_14237_));
 sky130_fd_sc_hd__and2b_1 _20963_ (.A_N(_14053_),
    .B(_14061_),
    .X(_14238_));
 sky130_fd_sc_hd__and2b_1 _20964_ (.A_N(_14052_),
    .B(_14062_),
    .X(_14239_));
 sky130_fd_sc_hd__and2b_1 _20965_ (.A_N(_14092_),
    .B(_14091_),
    .X(_14240_));
 sky130_fd_sc_hd__o21ba_1 _20966_ (.A1(_14054_),
    .A2(_14060_),
    .B1_N(_14057_),
    .X(_14241_));
 sky130_fd_sc_hd__o21ba_1 _20967_ (.A1(_14078_),
    .A2(_14082_),
    .B1_N(_14079_),
    .X(_14242_));
 sky130_fd_sc_hd__a22oi_1 _20968_ (.A1(_14055_),
    .A2(_14056_),
    .B1(_13446_),
    .B2(_11299_),
    .Y(_14243_));
 sky130_fd_sc_hd__and4_1 _20969_ (.A(_10783_),
    .B(_11201_),
    .C(_13285_),
    .D(_13445_),
    .X(_14244_));
 sky130_fd_sc_hd__nor2_1 _20970_ (.A(_14243_),
    .B(_14244_),
    .Y(_14245_));
 sky130_fd_sc_hd__nand2_1 _20971_ (.A(_11080_),
    .B(_13612_),
    .Y(_14246_));
 sky130_fd_sc_hd__xnor2_2 _20972_ (.A(_14245_),
    .B(_14246_),
    .Y(_14247_));
 sky130_fd_sc_hd__xnor2_1 _20973_ (.A(_14242_),
    .B(_14247_),
    .Y(_14248_));
 sky130_fd_sc_hd__xnor2_1 _20974_ (.A(_14241_),
    .B(_14248_),
    .Y(_14249_));
 sky130_fd_sc_hd__o21ai_1 _20975_ (.A1(_14240_),
    .A2(_14094_),
    .B1(_14249_),
    .Y(_14250_));
 sky130_fd_sc_hd__or3_1 _20976_ (.A(_14240_),
    .B(_14094_),
    .C(_14249_),
    .X(_14251_));
 sky130_fd_sc_hd__o211a_1 _20977_ (.A1(_14238_),
    .A2(_14239_),
    .B1(_14250_),
    .C1(_14251_),
    .X(_14252_));
 sky130_fd_sc_hd__a211oi_1 _20978_ (.A1(_14250_),
    .A2(_14251_),
    .B1(_14238_),
    .C1(_14239_),
    .Y(_14253_));
 sky130_fd_sc_hd__nor2_1 _20979_ (.A(_14252_),
    .B(_14253_),
    .Y(_14254_));
 sky130_fd_sc_hd__nor2_1 _20980_ (.A(_14064_),
    .B(_14066_),
    .Y(_14255_));
 sky130_fd_sc_hd__xnor2_2 _20981_ (.A(_14254_),
    .B(_14255_),
    .Y(_14256_));
 sky130_fd_sc_hd__xnor2_4 _20982_ (.A(_14237_),
    .B(_14256_),
    .Y(_14257_));
 sky130_fd_sc_hd__xnor2_2 _20983_ (.A(_14209_),
    .B(_14257_),
    .Y(_14258_));
 sky130_fd_sc_hd__xor2_4 _20984_ (.A(_14207_),
    .B(_14258_),
    .X(_14259_));
 sky130_fd_sc_hd__or2_2 _20985_ (.A(_14111_),
    .B(_14113_),
    .X(_14260_));
 sky130_fd_sc_hd__a21o_1 _20986_ (.A1(_14119_),
    .A2(_14141_),
    .B1(_14139_),
    .X(_14261_));
 sky130_fd_sc_hd__buf_2 _20987_ (.A(_13632_),
    .X(_14262_));
 sky130_fd_sc_hd__nand2_1 _20988_ (.A(_11138_),
    .B(_14262_),
    .Y(_14263_));
 sky130_fd_sc_hd__and4_1 _20989_ (.A(_13669_),
    .B(_11112_),
    .C(_13887_),
    .D(_12977_),
    .X(_14264_));
 sky130_fd_sc_hd__a22oi_1 _20990_ (.A1(_13665_),
    .A2(_14081_),
    .B1(_14077_),
    .B2(_13670_),
    .Y(_14265_));
 sky130_fd_sc_hd__nor2_1 _20991_ (.A(_14264_),
    .B(_14265_),
    .Y(_14266_));
 sky130_fd_sc_hd__xnor2_1 _20992_ (.A(_14263_),
    .B(_14266_),
    .Y(_14267_));
 sky130_fd_sc_hd__clkbuf_2 _20993_ (.A(_12983_),
    .X(_14268_));
 sky130_fd_sc_hd__buf_2 _20994_ (.A(_14268_),
    .X(_14269_));
 sky130_fd_sc_hd__nand2_1 _20995_ (.A(_11136_),
    .B(_14269_),
    .Y(_14270_));
 sky130_fd_sc_hd__and4_1 _20996_ (.A(_14086_),
    .B(_14087_),
    .C(_12145_),
    .D(_12274_),
    .X(_14271_));
 sky130_fd_sc_hd__clkbuf_2 _20997_ (.A(_12271_),
    .X(_14272_));
 sky130_fd_sc_hd__a22oi_2 _20998_ (.A1(_13900_),
    .A2(_13666_),
    .B1(_14272_),
    .B2(_13899_),
    .Y(_14273_));
 sky130_fd_sc_hd__nor2_1 _20999_ (.A(_14271_),
    .B(_14273_),
    .Y(_14274_));
 sky130_fd_sc_hd__xnor2_1 _21000_ (.A(_14270_),
    .B(_14274_),
    .Y(_14275_));
 sky130_fd_sc_hd__o21ba_1 _21001_ (.A1(_14085_),
    .A2(_14089_),
    .B1_N(_14088_),
    .X(_14276_));
 sky130_fd_sc_hd__xnor2_1 _21002_ (.A(_14275_),
    .B(_14276_),
    .Y(_14277_));
 sky130_fd_sc_hd__and2_1 _21003_ (.A(_14267_),
    .B(_14277_),
    .X(_14278_));
 sky130_fd_sc_hd__nor2_1 _21004_ (.A(_14267_),
    .B(_14277_),
    .Y(_14279_));
 sky130_fd_sc_hd__or2_2 _21005_ (.A(_14278_),
    .B(_14279_),
    .X(_14280_));
 sky130_fd_sc_hd__or2b_1 _21006_ (.A(_14101_),
    .B_N(_14108_),
    .X(_14281_));
 sky130_fd_sc_hd__nand2_1 _21007_ (.A(_14100_),
    .B(_14109_),
    .Y(_14282_));
 sky130_fd_sc_hd__clkbuf_4 _21008_ (.A(_11831_),
    .X(_14283_));
 sky130_fd_sc_hd__a31o_1 _21009_ (.A1(_11446_),
    .A2(_14283_),
    .A3(_14107_),
    .B1(_14104_),
    .X(_14284_));
 sky130_fd_sc_hd__o21ba_1 _21010_ (.A1(_14122_),
    .A2(_14125_),
    .B1_N(_14124_),
    .X(_14285_));
 sky130_fd_sc_hd__nand2_1 _21011_ (.A(_11560_),
    .B(_13674_),
    .Y(_14286_));
 sky130_fd_sc_hd__and4_1 _21012_ (.A(_14103_),
    .B(_13691_),
    .C(_11819_),
    .D(_11947_),
    .X(_14287_));
 sky130_fd_sc_hd__a22oi_1 _21013_ (.A1(_11927_),
    .A2(_11708_),
    .B1(_11831_),
    .B2(_14105_),
    .Y(_14288_));
 sky130_fd_sc_hd__nor2_1 _21014_ (.A(_14287_),
    .B(_14288_),
    .Y(_14289_));
 sky130_fd_sc_hd__xnor2_2 _21015_ (.A(_14286_),
    .B(_14289_),
    .Y(_14290_));
 sky130_fd_sc_hd__xnor2_1 _21016_ (.A(_14285_),
    .B(_14290_),
    .Y(_14291_));
 sky130_fd_sc_hd__xnor2_1 _21017_ (.A(_14284_),
    .B(_14291_),
    .Y(_14292_));
 sky130_fd_sc_hd__a21oi_1 _21018_ (.A1(_14281_),
    .A2(_14282_),
    .B1(_14292_),
    .Y(_14293_));
 sky130_fd_sc_hd__and3_1 _21019_ (.A(_14281_),
    .B(_14282_),
    .C(_14292_),
    .X(_14294_));
 sky130_fd_sc_hd__nor3_1 _21020_ (.A(_14280_),
    .B(_14293_),
    .C(_14294_),
    .Y(_14295_));
 sky130_fd_sc_hd__o21a_1 _21021_ (.A1(_14293_),
    .A2(_14294_),
    .B1(_14280_),
    .X(_14296_));
 sky130_fd_sc_hd__or2_2 _21022_ (.A(_14295_),
    .B(_14296_),
    .X(_14297_));
 sky130_fd_sc_hd__xnor2_2 _21023_ (.A(_14261_),
    .B(_14297_),
    .Y(_14298_));
 sky130_fd_sc_hd__xor2_4 _21024_ (.A(_14260_),
    .B(_14298_),
    .X(_14299_));
 sky130_fd_sc_hd__or2b_1 _21025_ (.A(_14136_),
    .B_N(_14135_),
    .X(_14300_));
 sky130_fd_sc_hd__a21bo_2 _21026_ (.A1(_14127_),
    .A2(_14137_),
    .B1_N(_14300_),
    .X(_14301_));
 sky130_fd_sc_hd__or3_1 _21027_ (.A(_14143_),
    .B(_14146_),
    .C(_14148_),
    .X(_14302_));
 sky130_fd_sc_hd__nand2_1 _21028_ (.A(_13690_),
    .B(_11771_),
    .Y(_14303_));
 sky130_fd_sc_hd__and4_1 _21029_ (.A(_11381_),
    .B(_11825_),
    .C(_14123_),
    .D(_13934_),
    .X(_14304_));
 sky130_fd_sc_hd__a22oi_2 _21030_ (.A1(_11491_),
    .A2(_11891_),
    .B1(_13937_),
    .B2(_11477_),
    .Y(_14305_));
 sky130_fd_sc_hd__nor2_1 _21031_ (.A(_14304_),
    .B(_14305_),
    .Y(_14306_));
 sky130_fd_sc_hd__xnor2_1 _21032_ (.A(_14303_),
    .B(_14306_),
    .Y(_14307_));
 sky130_fd_sc_hd__nand2_1 _21033_ (.A(_11278_),
    .B(_12227_),
    .Y(_14308_));
 sky130_fd_sc_hd__and4_1 _21034_ (.A(_11160_),
    .B(_11265_),
    .C(_12323_),
    .D(_13723_),
    .X(_14309_));
 sky130_fd_sc_hd__clkbuf_4 _21035_ (.A(_13376_),
    .X(_14310_));
 sky130_fd_sc_hd__a22oi_2 _21036_ (.A1(_11172_),
    .A2(_13942_),
    .B1(_14310_),
    .B2(_11056_),
    .Y(_14311_));
 sky130_fd_sc_hd__nor2_1 _21037_ (.A(_14309_),
    .B(_14311_),
    .Y(_14312_));
 sky130_fd_sc_hd__xnor2_1 _21038_ (.A(_14308_),
    .B(_14312_),
    .Y(_14313_));
 sky130_fd_sc_hd__o21ba_1 _21039_ (.A1(_14128_),
    .A2(_14133_),
    .B1_N(_14130_),
    .X(_14314_));
 sky130_fd_sc_hd__xnor2_1 _21040_ (.A(_14313_),
    .B(_14314_),
    .Y(_14315_));
 sky130_fd_sc_hd__xnor2_1 _21041_ (.A(_14307_),
    .B(_14315_),
    .Y(_14316_));
 sky130_fd_sc_hd__a21oi_1 _21042_ (.A1(_14302_),
    .A2(_14151_),
    .B1(_14316_),
    .Y(_14317_));
 sky130_fd_sc_hd__and3_1 _21043_ (.A(_14302_),
    .B(_14151_),
    .C(_14316_),
    .X(_14318_));
 sky130_fd_sc_hd__nor2_2 _21044_ (.A(_14317_),
    .B(_14318_),
    .Y(_14319_));
 sky130_fd_sc_hd__xor2_4 _21045_ (.A(_14301_),
    .B(_14319_),
    .X(_14320_));
 sky130_fd_sc_hd__o21ba_1 _21046_ (.A1(_14155_),
    .A2(_14157_),
    .B1_N(_14156_),
    .X(_14321_));
 sky130_fd_sc_hd__and4_2 _21047_ (.A(_11048_),
    .B(_10969_),
    .C(_13060_),
    .D(_13740_),
    .X(_14322_));
 sky130_fd_sc_hd__a22oi_2 _21048_ (.A1(_11280_),
    .A2(_12776_),
    .B1(_13960_),
    .B2(_11175_),
    .Y(_14323_));
 sky130_fd_sc_hd__clkbuf_2 _21049_ (.A(\genblk1.pcpi_mul.rs2[24] ),
    .X(_14324_));
 sky130_fd_sc_hd__and4bb_1 _21050_ (.A_N(_14322_),
    .B_N(_14323_),
    .C(_11043_),
    .D(_14324_),
    .X(_14325_));
 sky130_fd_sc_hd__o2bb2a_1 _21051_ (.A1_N(_11039_),
    .A2_N(_12585_),
    .B1(_14322_),
    .B2(_14323_),
    .X(_14326_));
 sky130_fd_sc_hd__nor2_1 _21052_ (.A(_14325_),
    .B(_14326_),
    .Y(_14327_));
 sky130_fd_sc_hd__xnor2_1 _21053_ (.A(_14321_),
    .B(_14327_),
    .Y(_14328_));
 sky130_fd_sc_hd__o21ai_2 _21054_ (.A1(_14144_),
    .A2(_14146_),
    .B1(_14328_),
    .Y(_14329_));
 sky130_fd_sc_hd__or3_1 _21055_ (.A(_14144_),
    .B(_14146_),
    .C(_14328_),
    .X(_14330_));
 sky130_fd_sc_hd__and2_2 _21056_ (.A(_14329_),
    .B(_14330_),
    .X(_14331_));
 sky130_fd_sc_hd__nand2_1 _21057_ (.A(_13959_),
    .B(_13055_),
    .Y(_14332_));
 sky130_fd_sc_hd__and4_1 _21058_ (.A(_11302_),
    .B(_11199_),
    .C(_13223_),
    .D(_13971_),
    .X(_14333_));
 sky130_fd_sc_hd__a22oi_2 _21059_ (.A1(_11404_),
    .A2(_13761_),
    .B1(_13972_),
    .B2(_11091_),
    .Y(_14334_));
 sky130_fd_sc_hd__nor2_1 _21060_ (.A(_14333_),
    .B(_14334_),
    .Y(_14335_));
 sky130_fd_sc_hd__xnor2_2 _21061_ (.A(_14332_),
    .B(_14335_),
    .Y(_14336_));
 sky130_fd_sc_hd__nand2_1 _21062_ (.A(_10666_),
    .B(_13541_),
    .Y(_14337_));
 sky130_fd_sc_hd__and2b_1 _21063_ (.A_N(_10754_),
    .B(_13802_),
    .X(_14338_));
 sky130_fd_sc_hd__nand2_1 _21064_ (.A(_10649_),
    .B(_13756_),
    .Y(_14339_));
 sky130_fd_sc_hd__xnor2_2 _21065_ (.A(_14338_),
    .B(_14339_),
    .Y(_14340_));
 sky130_fd_sc_hd__xnor2_2 _21066_ (.A(_14337_),
    .B(_14340_),
    .Y(_14341_));
 sky130_fd_sc_hd__clkbuf_2 _21067_ (.A(\genblk1.pcpi_mul.rs2[30] ),
    .X(_14342_));
 sky130_fd_sc_hd__buf_2 _21068_ (.A(_14342_),
    .X(_14343_));
 sky130_fd_sc_hd__and3_1 _21069_ (.A(_11778_),
    .B(_14168_),
    .C(_14162_),
    .X(_14344_));
 sky130_fd_sc_hd__a31o_1 _21070_ (.A1(_10676_),
    .A2(_14343_),
    .A3(_14164_),
    .B1(_14344_),
    .X(_14345_));
 sky130_fd_sc_hd__xor2_2 _21071_ (.A(_14341_),
    .B(_14345_),
    .X(_14346_));
 sky130_fd_sc_hd__xnor2_2 _21072_ (.A(_14336_),
    .B(_14346_),
    .Y(_14347_));
 sky130_fd_sc_hd__nand2_1 _21073_ (.A(_14165_),
    .B(_14170_),
    .Y(_14348_));
 sky130_fd_sc_hd__a21boi_2 _21074_ (.A1(_14159_),
    .A2(_14171_),
    .B1_N(_14348_),
    .Y(_14349_));
 sky130_fd_sc_hd__xnor2_2 _21075_ (.A(_14347_),
    .B(_14349_),
    .Y(_14350_));
 sky130_fd_sc_hd__xnor2_4 _21076_ (.A(_14331_),
    .B(_14350_),
    .Y(_14351_));
 sky130_fd_sc_hd__nand2_1 _21077_ (.A(_14172_),
    .B(_14174_),
    .Y(_14352_));
 sky130_fd_sc_hd__nor2_1 _21078_ (.A(_14172_),
    .B(_14174_),
    .Y(_14353_));
 sky130_fd_sc_hd__a21oi_2 _21079_ (.A1(_14153_),
    .A2(_14352_),
    .B1(_14353_),
    .Y(_14354_));
 sky130_fd_sc_hd__xnor2_4 _21080_ (.A(_14351_),
    .B(_14354_),
    .Y(_14355_));
 sky130_fd_sc_hd__xnor2_4 _21081_ (.A(_14320_),
    .B(_14355_),
    .Y(_14356_));
 sky130_fd_sc_hd__and2b_1 _21082_ (.A_N(_14178_),
    .B(_14176_),
    .X(_14357_));
 sky130_fd_sc_hd__a21oi_2 _21083_ (.A1(_14142_),
    .A2(_14179_),
    .B1(_14357_),
    .Y(_14358_));
 sky130_fd_sc_hd__xor2_4 _21084_ (.A(_14356_),
    .B(_14358_),
    .X(_14359_));
 sky130_fd_sc_hd__xor2_4 _21085_ (.A(_14299_),
    .B(_14359_),
    .X(_14360_));
 sky130_fd_sc_hd__nor2_1 _21086_ (.A(_14180_),
    .B(_14182_),
    .Y(_14361_));
 sky130_fd_sc_hd__a21oi_2 _21087_ (.A1(_14117_),
    .A2(_14183_),
    .B1(_14361_),
    .Y(_14362_));
 sky130_fd_sc_hd__xnor2_4 _21088_ (.A(_14360_),
    .B(_14362_),
    .Y(_14363_));
 sky130_fd_sc_hd__xnor2_4 _21089_ (.A(_14259_),
    .B(_14363_),
    .Y(_14364_));
 sky130_fd_sc_hd__nor2_1 _21090_ (.A(_14184_),
    .B(_14186_),
    .Y(_14365_));
 sky130_fd_sc_hd__a21oi_2 _21091_ (.A1(_14073_),
    .A2(_14187_),
    .B1(_14365_),
    .Y(_14366_));
 sky130_fd_sc_hd__xor2_4 _21092_ (.A(_14364_),
    .B(_14366_),
    .X(_14367_));
 sky130_fd_sc_hd__xnor2_4 _21093_ (.A(_14206_),
    .B(_14367_),
    .Y(_14368_));
 sky130_fd_sc_hd__nor2_1 _21094_ (.A(_14188_),
    .B(_14190_),
    .Y(_14369_));
 sky130_fd_sc_hd__a21oi_2 _21095_ (.A1(_14019_),
    .A2(_14191_),
    .B1(_14369_),
    .Y(_14370_));
 sky130_fd_sc_hd__xor2_4 _21096_ (.A(_14368_),
    .B(_14370_),
    .X(_14371_));
 sky130_fd_sc_hd__xnor2_4 _21097_ (.A(_14202_),
    .B(_14371_),
    .Y(_14372_));
 sky130_fd_sc_hd__and2b_1 _21098_ (.A_N(_14195_),
    .B(_14192_),
    .X(_14373_));
 sky130_fd_sc_hd__a21oi_4 _21099_ (.A1(_14015_),
    .A2(_14196_),
    .B1(_14373_),
    .Y(_14374_));
 sky130_fd_sc_hd__xnor2_4 _21100_ (.A(_14372_),
    .B(_14374_),
    .Y(_14375_));
 sky130_fd_sc_hd__and3b_1 _21101_ (.A_N(_14200_),
    .B(_14001_),
    .C(_14198_),
    .X(_14376_));
 sky130_fd_sc_hd__a21o_1 _21102_ (.A1(_14011_),
    .A2(_14198_),
    .B1(_14200_),
    .X(_14377_));
 sky130_fd_sc_hd__a21o_2 _21103_ (.A1(_14010_),
    .A2(_14376_),
    .B1(_14377_),
    .X(_14378_));
 sky130_fd_sc_hd__xnor2_4 _21104_ (.A(_14375_),
    .B(_14378_),
    .Y(_00080_));
 sky130_fd_sc_hd__nor2_1 _21105_ (.A(_14368_),
    .B(_14370_),
    .Y(_14379_));
 sky130_fd_sc_hd__a21oi_4 _21106_ (.A1(_14202_),
    .A2(_14371_),
    .B1(_14379_),
    .Y(_14380_));
 sky130_fd_sc_hd__o21a_2 _21107_ (.A1(_14042_),
    .A2(_14045_),
    .B1(_14204_),
    .X(_14381_));
 sky130_fd_sc_hd__and2b_1 _21108_ (.A_N(_14257_),
    .B(_14209_),
    .X(_14382_));
 sky130_fd_sc_hd__and2_1 _21109_ (.A(_14207_),
    .B(_14258_),
    .X(_14383_));
 sky130_fd_sc_hd__o21a_2 _21110_ (.A1(_14215_),
    .A2(_14236_),
    .B1(_14234_),
    .X(_14384_));
 sky130_fd_sc_hd__o21ba_2 _21111_ (.A1(_14382_),
    .A2(_14383_),
    .B1_N(_14384_),
    .X(_14385_));
 sky130_fd_sc_hd__or3b_1 _21112_ (.A(_14382_),
    .B(_14383_),
    .C_N(_14384_),
    .X(_14386_));
 sky130_fd_sc_hd__and2b_2 _21113_ (.A_N(_14385_),
    .B(_14386_),
    .X(_14387_));
 sky130_fd_sc_hd__nand2_1 _21114_ (.A(_14237_),
    .B(_14256_),
    .Y(_14388_));
 sky130_fd_sc_hd__o31a_2 _21115_ (.A1(_14252_),
    .A2(_14253_),
    .A3(_14255_),
    .B1(_14388_),
    .X(_14389_));
 sky130_fd_sc_hd__or2b_1 _21116_ (.A(_14297_),
    .B_N(_14261_),
    .X(_14390_));
 sky130_fd_sc_hd__a21bo_2 _21117_ (.A1(_14260_),
    .A2(_14298_),
    .B1_N(_14390_),
    .X(_14391_));
 sky130_fd_sc_hd__a31o_2 _21118_ (.A1(_11368_),
    .A2(_14214_),
    .A3(_14219_),
    .B1(_14025_),
    .X(_14392_));
 sky130_fd_sc_hd__nand2_1 _21119_ (.A(_14228_),
    .B(_14229_),
    .Y(_14393_));
 sky130_fd_sc_hd__nand2_2 _21120_ (.A(_10626_),
    .B(_14037_),
    .Y(_14394_));
 sky130_fd_sc_hd__xor2_4 _21121_ (.A(_14219_),
    .B(_14394_),
    .X(_14395_));
 sky130_vsdinv _21122_ (.A(_14395_),
    .Y(_14396_));
 sky130_fd_sc_hd__a22oi_1 _21123_ (.A1(_11385_),
    .A2(_14225_),
    .B1(_14210_),
    .B2(_11387_),
    .Y(_14397_));
 sky130_fd_sc_hd__buf_2 _21124_ (.A(\genblk1.pcpi_mul.rs1[31] ),
    .X(_14398_));
 sky130_fd_sc_hd__and4_1 _21125_ (.A(_10672_),
    .B(_11385_),
    .C(_13606_),
    .D(_14398_),
    .X(_14399_));
 sky130_fd_sc_hd__nor2_2 _21126_ (.A(_14397_),
    .B(_14399_),
    .Y(_14400_));
 sky130_fd_sc_hd__xnor2_1 _21127_ (.A(_14222_),
    .B(_14400_),
    .Y(_14401_));
 sky130_fd_sc_hd__o21ba_1 _21128_ (.A1(_14222_),
    .A2(_14224_),
    .B1_N(_14226_),
    .X(_14402_));
 sky130_fd_sc_hd__xnor2_1 _21129_ (.A(_14401_),
    .B(_14402_),
    .Y(_14403_));
 sky130_fd_sc_hd__nand2_1 _21130_ (.A(_14396_),
    .B(_14403_),
    .Y(_14404_));
 sky130_fd_sc_hd__or2_1 _21131_ (.A(_14396_),
    .B(_14403_),
    .X(_14405_));
 sky130_fd_sc_hd__nand2_1 _21132_ (.A(_14404_),
    .B(_14405_),
    .Y(_14406_));
 sky130_fd_sc_hd__a21oi_1 _21133_ (.A1(_14393_),
    .A2(_14231_),
    .B1(_14406_),
    .Y(_14407_));
 sky130_fd_sc_hd__nand3_1 _21134_ (.A(_14393_),
    .B(_14231_),
    .C(_14406_),
    .Y(_14408_));
 sky130_fd_sc_hd__or2b_1 _21135_ (.A(_14407_),
    .B_N(_14408_),
    .X(_14409_));
 sky130_fd_sc_hd__xnor2_2 _21136_ (.A(_14392_),
    .B(_14409_),
    .Y(_14410_));
 sky130_fd_sc_hd__and2b_1 _21137_ (.A_N(_14242_),
    .B(_14247_),
    .X(_14411_));
 sky130_fd_sc_hd__and2b_1 _21138_ (.A_N(_14241_),
    .B(_14248_),
    .X(_14412_));
 sky130_fd_sc_hd__and2b_1 _21139_ (.A_N(_14276_),
    .B(_14275_),
    .X(_14413_));
 sky130_fd_sc_hd__o21ba_1 _21140_ (.A1(_14243_),
    .A2(_14246_),
    .B1_N(_14244_),
    .X(_14414_));
 sky130_fd_sc_hd__o21ba_1 _21141_ (.A1(_14263_),
    .A2(_14265_),
    .B1_N(_14264_),
    .X(_14415_));
 sky130_fd_sc_hd__a22oi_1 _21142_ (.A1(_14055_),
    .A2(_13838_),
    .B1(_13839_),
    .B2(_13863_),
    .Y(_14416_));
 sky130_fd_sc_hd__clkbuf_2 _21143_ (.A(_12980_),
    .X(_14417_));
 sky130_fd_sc_hd__clkbuf_2 _21144_ (.A(_13128_),
    .X(_14418_));
 sky130_fd_sc_hd__and4_1 _21145_ (.A(_11299_),
    .B(_11197_),
    .C(_14417_),
    .D(_14418_),
    .X(_14419_));
 sky130_fd_sc_hd__nor2_1 _21146_ (.A(_14416_),
    .B(_14419_),
    .Y(_14420_));
 sky130_fd_sc_hd__nand2_1 _21147_ (.A(_11080_),
    .B(_13814_),
    .Y(_14421_));
 sky130_fd_sc_hd__xnor2_1 _21148_ (.A(_14420_),
    .B(_14421_),
    .Y(_14422_));
 sky130_fd_sc_hd__xnor2_1 _21149_ (.A(_14415_),
    .B(_14422_),
    .Y(_14423_));
 sky130_fd_sc_hd__xnor2_1 _21150_ (.A(_14414_),
    .B(_14423_),
    .Y(_14424_));
 sky130_fd_sc_hd__o21ai_1 _21151_ (.A1(_14413_),
    .A2(_14278_),
    .B1(_14424_),
    .Y(_14425_));
 sky130_fd_sc_hd__or3_1 _21152_ (.A(_14413_),
    .B(_14278_),
    .C(_14424_),
    .X(_14426_));
 sky130_fd_sc_hd__o211a_1 _21153_ (.A1(_14411_),
    .A2(_14412_),
    .B1(_14425_),
    .C1(_14426_),
    .X(_14427_));
 sky130_fd_sc_hd__a211oi_1 _21154_ (.A1(_14425_),
    .A2(_14426_),
    .B1(_14411_),
    .C1(_14412_),
    .Y(_14428_));
 sky130_fd_sc_hd__nor2_1 _21155_ (.A(_14427_),
    .B(_14428_),
    .Y(_14429_));
 sky130_vsdinv _21156_ (.A(_14250_),
    .Y(_14430_));
 sky130_fd_sc_hd__nor2_1 _21157_ (.A(_14430_),
    .B(_14252_),
    .Y(_14431_));
 sky130_fd_sc_hd__xnor2_2 _21158_ (.A(_14429_),
    .B(_14431_),
    .Y(_14432_));
 sky130_fd_sc_hd__xnor2_2 _21159_ (.A(_14410_),
    .B(_14432_),
    .Y(_14433_));
 sky130_fd_sc_hd__xnor2_2 _21160_ (.A(_14391_),
    .B(_14433_),
    .Y(_14434_));
 sky130_fd_sc_hd__xnor2_4 _21161_ (.A(_14389_),
    .B(_14434_),
    .Y(_14435_));
 sky130_fd_sc_hd__or2_2 _21162_ (.A(_14293_),
    .B(_14295_),
    .X(_14436_));
 sky130_fd_sc_hd__a21o_1 _21163_ (.A1(_14301_),
    .A2(_14319_),
    .B1(_14317_),
    .X(_14437_));
 sky130_fd_sc_hd__buf_2 _21164_ (.A(_14056_),
    .X(_14438_));
 sky130_fd_sc_hd__nand2_1 _21165_ (.A(_11138_),
    .B(_14438_),
    .Y(_14439_));
 sky130_fd_sc_hd__and4_1 _21166_ (.A(_13661_),
    .B(_13662_),
    .C(_12977_),
    .D(_13864_),
    .X(_14440_));
 sky130_fd_sc_hd__a22oi_2 _21167_ (.A1(_11109_),
    .A2(_14077_),
    .B1(_14262_),
    .B2(_10958_),
    .Y(_14441_));
 sky130_fd_sc_hd__nor2_1 _21168_ (.A(_14440_),
    .B(_14441_),
    .Y(_14442_));
 sky130_fd_sc_hd__xnor2_1 _21169_ (.A(_14439_),
    .B(_14442_),
    .Y(_14443_));
 sky130_fd_sc_hd__clkbuf_4 _21170_ (.A(_12416_),
    .X(_14444_));
 sky130_fd_sc_hd__nand2_1 _21171_ (.A(_11136_),
    .B(_14444_),
    .Y(_14445_));
 sky130_fd_sc_hd__and4_1 _21172_ (.A(_14086_),
    .B(_14087_),
    .C(_12274_),
    .D(_14268_),
    .X(_14446_));
 sky130_fd_sc_hd__a22oi_2 _21173_ (.A1(_13900_),
    .A2(_14272_),
    .B1(_13890_),
    .B2(_13899_),
    .Y(_14447_));
 sky130_fd_sc_hd__nor2_1 _21174_ (.A(_14446_),
    .B(_14447_),
    .Y(_14448_));
 sky130_fd_sc_hd__xnor2_1 _21175_ (.A(_14445_),
    .B(_14448_),
    .Y(_14449_));
 sky130_fd_sc_hd__o21ba_1 _21176_ (.A1(_14270_),
    .A2(_14273_),
    .B1_N(_14271_),
    .X(_14450_));
 sky130_fd_sc_hd__xnor2_1 _21177_ (.A(_14449_),
    .B(_14450_),
    .Y(_14451_));
 sky130_fd_sc_hd__and2_1 _21178_ (.A(_14443_),
    .B(_14451_),
    .X(_14452_));
 sky130_fd_sc_hd__nor2_1 _21179_ (.A(_14443_),
    .B(_14451_),
    .Y(_14453_));
 sky130_fd_sc_hd__or2_2 _21180_ (.A(_14452_),
    .B(_14453_),
    .X(_14454_));
 sky130_fd_sc_hd__or2b_1 _21181_ (.A(_14285_),
    .B_N(_14290_),
    .X(_14455_));
 sky130_fd_sc_hd__nand2_1 _21182_ (.A(_14284_),
    .B(_14291_),
    .Y(_14456_));
 sky130_fd_sc_hd__buf_2 _21183_ (.A(_11959_),
    .X(_14457_));
 sky130_fd_sc_hd__a31o_2 _21184_ (.A1(_11446_),
    .A2(_14457_),
    .A3(_14289_),
    .B1(_14287_),
    .X(_14458_));
 sky130_fd_sc_hd__o21ba_1 _21185_ (.A1(_14303_),
    .A2(_14305_),
    .B1_N(_14304_),
    .X(_14459_));
 sky130_fd_sc_hd__nand2_1 _21186_ (.A(_11775_),
    .B(_12413_),
    .Y(_14460_));
 sky130_fd_sc_hd__and4_1 _21187_ (.A(_14103_),
    .B(_13691_),
    .C(_11947_),
    .D(_12070_),
    .X(_14461_));
 sky130_fd_sc_hd__a22oi_1 _21188_ (.A1(_11927_),
    .A2(_13679_),
    .B1(_13901_),
    .B2(_14105_),
    .Y(_14462_));
 sky130_fd_sc_hd__nor2_1 _21189_ (.A(_14461_),
    .B(_14462_),
    .Y(_14463_));
 sky130_fd_sc_hd__xnor2_2 _21190_ (.A(_14460_),
    .B(_14463_),
    .Y(_14464_));
 sky130_fd_sc_hd__xnor2_1 _21191_ (.A(_14459_),
    .B(_14464_),
    .Y(_14465_));
 sky130_fd_sc_hd__xnor2_1 _21192_ (.A(_14458_),
    .B(_14465_),
    .Y(_14466_));
 sky130_fd_sc_hd__a21oi_1 _21193_ (.A1(_14455_),
    .A2(_14456_),
    .B1(_14466_),
    .Y(_14467_));
 sky130_fd_sc_hd__and3_1 _21194_ (.A(_14455_),
    .B(_14456_),
    .C(_14466_),
    .X(_14468_));
 sky130_fd_sc_hd__nor3_1 _21195_ (.A(_14454_),
    .B(_14467_),
    .C(_14468_),
    .Y(_14469_));
 sky130_fd_sc_hd__o21a_1 _21196_ (.A1(_14467_),
    .A2(_14468_),
    .B1(_14454_),
    .X(_14470_));
 sky130_fd_sc_hd__or2_1 _21197_ (.A(_14469_),
    .B(_14470_),
    .X(_14471_));
 sky130_fd_sc_hd__xnor2_2 _21198_ (.A(_14437_),
    .B(_14471_),
    .Y(_14472_));
 sky130_fd_sc_hd__xor2_4 _21199_ (.A(_14436_),
    .B(_14472_),
    .X(_14473_));
 sky130_fd_sc_hd__or2b_1 _21200_ (.A(_14314_),
    .B_N(_14313_),
    .X(_14474_));
 sky130_fd_sc_hd__nand2_1 _21201_ (.A(_14307_),
    .B(_14315_),
    .Y(_14475_));
 sky130_fd_sc_hd__or3_2 _21202_ (.A(_14321_),
    .B(_14325_),
    .C(_14326_),
    .X(_14476_));
 sky130_fd_sc_hd__nand2_1 _21203_ (.A(_13919_),
    .B(_13711_),
    .Y(_14477_));
 sky130_fd_sc_hd__and4_1 _21204_ (.A(_11591_),
    .B(_13695_),
    .C(_11896_),
    .D(_13934_),
    .X(_14478_));
 sky130_fd_sc_hd__a22oi_2 _21205_ (.A1(_13690_),
    .A2(_13936_),
    .B1(_13937_),
    .B2(_11826_),
    .Y(_14479_));
 sky130_fd_sc_hd__nor2_1 _21206_ (.A(_14478_),
    .B(_14479_),
    .Y(_14480_));
 sky130_fd_sc_hd__xnor2_1 _21207_ (.A(_14477_),
    .B(_14480_),
    .Y(_14481_));
 sky130_fd_sc_hd__buf_2 _21208_ (.A(_12226_),
    .X(_14482_));
 sky130_fd_sc_hd__nand2_1 _21209_ (.A(_11477_),
    .B(_14482_),
    .Y(_14483_));
 sky130_fd_sc_hd__and4_1 _21210_ (.A(_11601_),
    .B(_11372_),
    .C(_14131_),
    .D(_13374_),
    .X(_14484_));
 sky130_fd_sc_hd__a22oi_2 _21211_ (.A1(_12343_),
    .A2(_12323_),
    .B1(_14129_),
    .B2(_11265_),
    .Y(_14485_));
 sky130_fd_sc_hd__nor2_1 _21212_ (.A(_14484_),
    .B(_14485_),
    .Y(_14486_));
 sky130_fd_sc_hd__xnor2_1 _21213_ (.A(_14483_),
    .B(_14486_),
    .Y(_14487_));
 sky130_fd_sc_hd__o21ba_1 _21214_ (.A1(_14308_),
    .A2(_14311_),
    .B1_N(_14309_),
    .X(_14488_));
 sky130_fd_sc_hd__xnor2_1 _21215_ (.A(_14487_),
    .B(_14488_),
    .Y(_14489_));
 sky130_fd_sc_hd__xnor2_1 _21216_ (.A(_14481_),
    .B(_14489_),
    .Y(_14490_));
 sky130_fd_sc_hd__a21oi_1 _21217_ (.A1(_14476_),
    .A2(_14329_),
    .B1(_14490_),
    .Y(_14491_));
 sky130_fd_sc_hd__and3_1 _21218_ (.A(_14476_),
    .B(_14329_),
    .C(_14490_),
    .X(_14492_));
 sky130_fd_sc_hd__a211o_1 _21219_ (.A1(_14474_),
    .A2(_14475_),
    .B1(_14491_),
    .C1(_14492_),
    .X(_14493_));
 sky130_fd_sc_hd__o211ai_1 _21220_ (.A1(_14491_),
    .A2(_14492_),
    .B1(_14474_),
    .C1(_14475_),
    .Y(_14494_));
 sky130_fd_sc_hd__and2_2 _21221_ (.A(_14493_),
    .B(_14494_),
    .X(_14495_));
 sky130_fd_sc_hd__o21ba_1 _21222_ (.A1(_14332_),
    .A2(_14334_),
    .B1_N(_14333_),
    .X(_14496_));
 sky130_fd_sc_hd__and4_2 _21223_ (.A(_11036_),
    .B(_11038_),
    .C(_13558_),
    .D(_13740_),
    .X(_14497_));
 sky130_fd_sc_hd__a22oi_2 _21224_ (.A1(_11269_),
    .A2(_12771_),
    .B1(_13960_),
    .B2(_11280_),
    .Y(_14498_));
 sky130_fd_sc_hd__clkbuf_2 _21225_ (.A(_12775_),
    .X(_14499_));
 sky130_fd_sc_hd__and4bb_1 _21226_ (.A_N(_14497_),
    .B_N(_14498_),
    .C(_11728_),
    .D(_14499_),
    .X(_14500_));
 sky130_fd_sc_hd__o2bb2a_1 _21227_ (.A1_N(_11068_),
    .A2_N(_12585_),
    .B1(_14497_),
    .B2(_14498_),
    .X(_14501_));
 sky130_fd_sc_hd__nor2_1 _21228_ (.A(_14500_),
    .B(_14501_),
    .Y(_14502_));
 sky130_fd_sc_hd__xnor2_1 _21229_ (.A(_14496_),
    .B(_14502_),
    .Y(_14503_));
 sky130_fd_sc_hd__o21ai_2 _21230_ (.A1(_14322_),
    .A2(_14325_),
    .B1(_14503_),
    .Y(_14504_));
 sky130_fd_sc_hd__or3_1 _21231_ (.A(_14322_),
    .B(_14325_),
    .C(_14503_),
    .X(_14505_));
 sky130_fd_sc_hd__and2_2 _21232_ (.A(_14504_),
    .B(_14505_),
    .X(_14506_));
 sky130_fd_sc_hd__nand2_1 _21233_ (.A(_11050_),
    .B(_13226_),
    .Y(_14507_));
 sky130_fd_sc_hd__clkbuf_2 _21234_ (.A(_13545_),
    .X(_14508_));
 sky130_fd_sc_hd__and4_1 _21235_ (.A(_11193_),
    .B(_11405_),
    .C(_13761_),
    .D(_14508_),
    .X(_14509_));
 sky130_fd_sc_hd__clkbuf_4 _21236_ (.A(_13765_),
    .X(_14510_));
 sky130_fd_sc_hd__a22oi_2 _21237_ (.A1(_13959_),
    .A2(_13970_),
    .B1(_14510_),
    .B2(_12361_),
    .Y(_14511_));
 sky130_fd_sc_hd__nor2_1 _21238_ (.A(_14509_),
    .B(_14511_),
    .Y(_14512_));
 sky130_fd_sc_hd__xnor2_2 _21239_ (.A(_14507_),
    .B(_14512_),
    .Y(_14513_));
 sky130_fd_sc_hd__nand2_1 _21240_ (.A(_11091_),
    .B(_13541_),
    .Y(_14514_));
 sky130_fd_sc_hd__and2b_1 _21241_ (.A_N(_10717_),
    .B(_13802_),
    .X(_14515_));
 sky130_fd_sc_hd__nand2_1 _21242_ (.A(_10742_),
    .B(_13756_),
    .Y(_14516_));
 sky130_fd_sc_hd__xnor2_2 _21243_ (.A(_14515_),
    .B(_14516_),
    .Y(_14517_));
 sky130_fd_sc_hd__xnor2_2 _21244_ (.A(_14514_),
    .B(_14517_),
    .Y(_14518_));
 sky130_fd_sc_hd__and3_1 _21245_ (.A(_10650_),
    .B(_14168_),
    .C(_14338_),
    .X(_14519_));
 sky130_fd_sc_hd__a31o_1 _21246_ (.A1(_11245_),
    .A2(_14343_),
    .A3(_14340_),
    .B1(_14519_),
    .X(_14520_));
 sky130_fd_sc_hd__xor2_2 _21247_ (.A(_14518_),
    .B(_14520_),
    .X(_14521_));
 sky130_fd_sc_hd__xnor2_2 _21248_ (.A(_14513_),
    .B(_14521_),
    .Y(_14522_));
 sky130_fd_sc_hd__nand2_1 _21249_ (.A(_14341_),
    .B(_14345_),
    .Y(_14523_));
 sky130_fd_sc_hd__a21boi_2 _21250_ (.A1(_14336_),
    .A2(_14346_),
    .B1_N(_14523_),
    .Y(_14524_));
 sky130_fd_sc_hd__xnor2_2 _21251_ (.A(_14522_),
    .B(_14524_),
    .Y(_14525_));
 sky130_fd_sc_hd__xnor2_4 _21252_ (.A(_14506_),
    .B(_14525_),
    .Y(_14526_));
 sky130_fd_sc_hd__nand2_1 _21253_ (.A(_14347_),
    .B(_14349_),
    .Y(_14527_));
 sky130_fd_sc_hd__nor2_1 _21254_ (.A(_14347_),
    .B(_14349_),
    .Y(_14528_));
 sky130_fd_sc_hd__a21oi_2 _21255_ (.A1(_14331_),
    .A2(_14527_),
    .B1(_14528_),
    .Y(_14529_));
 sky130_fd_sc_hd__xnor2_4 _21256_ (.A(_14526_),
    .B(_14529_),
    .Y(_14530_));
 sky130_fd_sc_hd__xnor2_4 _21257_ (.A(_14495_),
    .B(_14530_),
    .Y(_14531_));
 sky130_fd_sc_hd__and2b_1 _21258_ (.A_N(_14354_),
    .B(_14351_),
    .X(_14532_));
 sky130_fd_sc_hd__a21oi_2 _21259_ (.A1(_14320_),
    .A2(_14355_),
    .B1(_14532_),
    .Y(_14533_));
 sky130_fd_sc_hd__xor2_4 _21260_ (.A(_14531_),
    .B(_14533_),
    .X(_14534_));
 sky130_fd_sc_hd__xor2_4 _21261_ (.A(_14473_),
    .B(_14534_),
    .X(_14535_));
 sky130_fd_sc_hd__nor2_1 _21262_ (.A(_14356_),
    .B(_14358_),
    .Y(_14536_));
 sky130_fd_sc_hd__a21oi_2 _21263_ (.A1(_14299_),
    .A2(_14359_),
    .B1(_14536_),
    .Y(_14537_));
 sky130_fd_sc_hd__xnor2_4 _21264_ (.A(_14535_),
    .B(_14537_),
    .Y(_14538_));
 sky130_fd_sc_hd__xnor2_4 _21265_ (.A(_14435_),
    .B(_14538_),
    .Y(_14539_));
 sky130_fd_sc_hd__or2b_1 _21266_ (.A(_14362_),
    .B_N(_14360_),
    .X(_14540_));
 sky130_fd_sc_hd__a21boi_4 _21267_ (.A1(_14259_),
    .A2(_14363_),
    .B1_N(_14540_),
    .Y(_14541_));
 sky130_fd_sc_hd__xor2_4 _21268_ (.A(_14539_),
    .B(_14541_),
    .X(_14542_));
 sky130_fd_sc_hd__xnor2_4 _21269_ (.A(_14387_),
    .B(_14542_),
    .Y(_14543_));
 sky130_fd_sc_hd__nor2_1 _21270_ (.A(_14364_),
    .B(_14366_),
    .Y(_14544_));
 sky130_fd_sc_hd__a21oi_2 _21271_ (.A1(_14206_),
    .A2(_14367_),
    .B1(_14544_),
    .Y(_14545_));
 sky130_fd_sc_hd__xor2_4 _21272_ (.A(_14543_),
    .B(_14545_),
    .X(_14546_));
 sky130_fd_sc_hd__xnor2_4 _21273_ (.A(_14381_),
    .B(_14546_),
    .Y(_14547_));
 sky130_fd_sc_hd__xor2_4 _21274_ (.A(_14380_),
    .B(_14547_),
    .X(_14548_));
 sky130_fd_sc_hd__nand2_1 _21275_ (.A(_14372_),
    .B(_14374_),
    .Y(_14549_));
 sky130_fd_sc_hd__nor2_1 _21276_ (.A(_14372_),
    .B(_14374_),
    .Y(_14550_));
 sky130_fd_sc_hd__a21oi_2 _21277_ (.A1(_14549_),
    .A2(_14378_),
    .B1(_14550_),
    .Y(_14551_));
 sky130_fd_sc_hd__xnor2_4 _21278_ (.A(_14548_),
    .B(_14551_),
    .Y(_00081_));
 sky130_fd_sc_hd__or2b_1 _21279_ (.A(_14433_),
    .B_N(_14391_),
    .X(_14552_));
 sky130_fd_sc_hd__or2b_1 _21280_ (.A(_14389_),
    .B_N(_14434_),
    .X(_14553_));
 sky130_fd_sc_hd__a21oi_1 _21281_ (.A1(_14392_),
    .A2(_14408_),
    .B1(_14407_),
    .Y(_14554_));
 sky130_fd_sc_hd__a21oi_2 _21282_ (.A1(_14552_),
    .A2(_14553_),
    .B1(_14554_),
    .Y(_14555_));
 sky130_fd_sc_hd__and3_1 _21283_ (.A(_14552_),
    .B(_14553_),
    .C(_14554_),
    .X(_14556_));
 sky130_fd_sc_hd__nor2_1 _21284_ (.A(_14555_),
    .B(_14556_),
    .Y(_14557_));
 sky130_fd_sc_hd__and2b_1 _21285_ (.A_N(_14431_),
    .B(_14429_),
    .X(_14558_));
 sky130_fd_sc_hd__a21oi_2 _21286_ (.A1(_14410_),
    .A2(_14432_),
    .B1(_14558_),
    .Y(_14559_));
 sky130_fd_sc_hd__or2b_1 _21287_ (.A(_14471_),
    .B_N(_14437_),
    .X(_14560_));
 sky130_fd_sc_hd__a21bo_1 _21288_ (.A1(_14436_),
    .A2(_14472_),
    .B1_N(_14560_),
    .X(_14561_));
 sky130_fd_sc_hd__clkbuf_4 _21289_ (.A(_14026_),
    .X(_14562_));
 sky130_fd_sc_hd__clkbuf_2 _21290_ (.A(_14562_),
    .X(_14563_));
 sky130_fd_sc_hd__buf_2 _21291_ (.A(_14563_),
    .X(_14564_));
 sky130_fd_sc_hd__clkbuf_4 _21292_ (.A(_14564_),
    .X(_14565_));
 sky130_fd_sc_hd__a31o_2 _21293_ (.A1(_11368_),
    .A2(_14565_),
    .A3(_14219_),
    .B1(_14025_),
    .X(_14566_));
 sky130_fd_sc_hd__clkbuf_4 _21294_ (.A(_14566_),
    .X(_14567_));
 sky130_fd_sc_hd__or2b_1 _21295_ (.A(_14402_),
    .B_N(_14401_),
    .X(_14568_));
 sky130_fd_sc_hd__a31o_1 _21296_ (.A1(_10585_),
    .A2(_14038_),
    .A3(_14400_),
    .B1(_14399_),
    .X(_14569_));
 sky130_fd_sc_hd__clkbuf_4 _21297_ (.A(_14024_),
    .X(_14570_));
 sky130_fd_sc_hd__a22o_1 _21298_ (.A1(_14223_),
    .A2(_13827_),
    .B1(_14570_),
    .B2(_11387_),
    .X(_14571_));
 sky130_fd_sc_hd__nand4_1 _21299_ (.A(_10663_),
    .B(_14223_),
    .C(_13827_),
    .D(_14037_),
    .Y(_01500_));
 sky130_fd_sc_hd__nand2_1 _21300_ (.A(_14571_),
    .B(_01500_),
    .Y(_01501_));
 sky130_fd_sc_hd__xor2_1 _21301_ (.A(_14222_),
    .B(_01501_),
    .X(_01502_));
 sky130_fd_sc_hd__xnor2_1 _21302_ (.A(_14569_),
    .B(_01502_),
    .Y(_01503_));
 sky130_fd_sc_hd__or2_1 _21303_ (.A(_14395_),
    .B(_01503_),
    .X(_01504_));
 sky130_fd_sc_hd__nand2_1 _21304_ (.A(_14395_),
    .B(_01503_),
    .Y(_01505_));
 sky130_fd_sc_hd__nand2_1 _21305_ (.A(_01504_),
    .B(_01505_),
    .Y(_01506_));
 sky130_fd_sc_hd__a21oi_1 _21306_ (.A1(_14568_),
    .A2(_14404_),
    .B1(_01506_),
    .Y(_01507_));
 sky130_fd_sc_hd__and3_1 _21307_ (.A(_14568_),
    .B(_14404_),
    .C(_01506_),
    .X(_01508_));
 sky130_fd_sc_hd__nor2_1 _21308_ (.A(_01507_),
    .B(_01508_),
    .Y(_01509_));
 sky130_fd_sc_hd__xnor2_1 _21309_ (.A(_14567_),
    .B(_01509_),
    .Y(_01510_));
 sky130_fd_sc_hd__or2b_1 _21310_ (.A(_14415_),
    .B_N(_14422_),
    .X(_01511_));
 sky130_fd_sc_hd__or2b_1 _21311_ (.A(_14414_),
    .B_N(_14423_),
    .X(_01512_));
 sky130_fd_sc_hd__and2b_1 _21312_ (.A_N(_14450_),
    .B(_14449_),
    .X(_01513_));
 sky130_fd_sc_hd__o21ba_1 _21313_ (.A1(_14416_),
    .A2(_14421_),
    .B1_N(_14419_),
    .X(_01514_));
 sky130_fd_sc_hd__o21ba_1 _21314_ (.A1(_14439_),
    .A2(_14441_),
    .B1_N(_14440_),
    .X(_01515_));
 sky130_fd_sc_hd__clkbuf_2 _21315_ (.A(_13281_),
    .X(_01516_));
 sky130_fd_sc_hd__a22oi_1 _21316_ (.A1(_14055_),
    .A2(_01516_),
    .B1(_14033_),
    .B2(_13863_),
    .Y(_01517_));
 sky130_fd_sc_hd__and4_1 _21317_ (.A(_11299_),
    .B(_11197_),
    .C(_14418_),
    .D(_13813_),
    .X(_01518_));
 sky130_fd_sc_hd__nor2_1 _21318_ (.A(_01517_),
    .B(_01518_),
    .Y(_01519_));
 sky130_fd_sc_hd__nand2_1 _21319_ (.A(_11080_),
    .B(_13829_),
    .Y(_01520_));
 sky130_fd_sc_hd__xnor2_2 _21320_ (.A(_01519_),
    .B(_01520_),
    .Y(_01521_));
 sky130_fd_sc_hd__xnor2_1 _21321_ (.A(_01515_),
    .B(_01521_),
    .Y(_01522_));
 sky130_fd_sc_hd__xnor2_1 _21322_ (.A(_01514_),
    .B(_01522_),
    .Y(_01523_));
 sky130_fd_sc_hd__o21a_1 _21323_ (.A1(_01513_),
    .A2(_14452_),
    .B1(_01523_),
    .X(_01524_));
 sky130_fd_sc_hd__nor3_1 _21324_ (.A(_01513_),
    .B(_14452_),
    .C(_01523_),
    .Y(_01525_));
 sky130_fd_sc_hd__a211oi_2 _21325_ (.A1(_01511_),
    .A2(_01512_),
    .B1(_01524_),
    .C1(_01525_),
    .Y(_01526_));
 sky130_fd_sc_hd__o211a_1 _21326_ (.A1(_01524_),
    .A2(_01525_),
    .B1(_01511_),
    .C1(_01512_),
    .X(_01527_));
 sky130_fd_sc_hd__or2_1 _21327_ (.A(_01526_),
    .B(_01527_),
    .X(_01528_));
 sky130_vsdinv _21328_ (.A(_14425_),
    .Y(_01529_));
 sky130_fd_sc_hd__nor2_1 _21329_ (.A(_01529_),
    .B(_14427_),
    .Y(_01530_));
 sky130_fd_sc_hd__xnor2_1 _21330_ (.A(_01528_),
    .B(_01530_),
    .Y(_01531_));
 sky130_fd_sc_hd__xnor2_1 _21331_ (.A(_01510_),
    .B(_01531_),
    .Y(_01532_));
 sky130_fd_sc_hd__xnor2_1 _21332_ (.A(_14561_),
    .B(_01532_),
    .Y(_01533_));
 sky130_fd_sc_hd__xnor2_2 _21333_ (.A(_14559_),
    .B(_01533_),
    .Y(_01534_));
 sky130_fd_sc_hd__nor2_1 _21334_ (.A(_14467_),
    .B(_14469_),
    .Y(_01535_));
 sky130_fd_sc_hd__a21o_1 _21335_ (.A1(_14476_),
    .A2(_14329_),
    .B1(_14490_),
    .X(_01536_));
 sky130_fd_sc_hd__nand2_1 _21336_ (.A(_10894_),
    .B(_14059_),
    .Y(_01537_));
 sky130_fd_sc_hd__buf_2 _21337_ (.A(_14056_),
    .X(_01538_));
 sky130_fd_sc_hd__and4_1 _21338_ (.A(_10958_),
    .B(_13665_),
    .C(_13861_),
    .D(_01538_),
    .X(_01539_));
 sky130_fd_sc_hd__clkbuf_2 _21339_ (.A(_13637_),
    .X(_01540_));
 sky130_fd_sc_hd__a22oi_1 _21340_ (.A1(_11109_),
    .A2(_01540_),
    .B1(_14438_),
    .B2(_10958_),
    .Y(_01541_));
 sky130_fd_sc_hd__nor2_1 _21341_ (.A(_01539_),
    .B(_01541_),
    .Y(_01542_));
 sky130_fd_sc_hd__xnor2_2 _21342_ (.A(_01537_),
    .B(_01542_),
    .Y(_01543_));
 sky130_fd_sc_hd__clkbuf_4 _21343_ (.A(_12977_),
    .X(_01544_));
 sky130_fd_sc_hd__nand2_1 _21344_ (.A(_11233_),
    .B(_01544_),
    .Y(_01545_));
 sky130_fd_sc_hd__and4_1 _21345_ (.A(_11242_),
    .B(_13903_),
    .C(_12694_),
    .D(_13887_),
    .X(_01546_));
 sky130_fd_sc_hd__buf_4 _21346_ (.A(_14087_),
    .X(_01547_));
 sky130_fd_sc_hd__a22oi_1 _21347_ (.A1(_01547_),
    .A2(_14269_),
    .B1(_14081_),
    .B2(_11237_),
    .Y(_01548_));
 sky130_fd_sc_hd__nor2_1 _21348_ (.A(_01546_),
    .B(_01548_),
    .Y(_01549_));
 sky130_fd_sc_hd__xnor2_1 _21349_ (.A(_01545_),
    .B(_01549_),
    .Y(_01550_));
 sky130_fd_sc_hd__o21ba_1 _21350_ (.A1(_14445_),
    .A2(_14447_),
    .B1_N(_14446_),
    .X(_01551_));
 sky130_fd_sc_hd__xnor2_1 _21351_ (.A(_01550_),
    .B(_01551_),
    .Y(_01552_));
 sky130_fd_sc_hd__and2_1 _21352_ (.A(_01543_),
    .B(_01552_),
    .X(_01553_));
 sky130_fd_sc_hd__nor2_1 _21353_ (.A(_01543_),
    .B(_01552_),
    .Y(_01554_));
 sky130_fd_sc_hd__or2_2 _21354_ (.A(_01553_),
    .B(_01554_),
    .X(_01555_));
 sky130_fd_sc_hd__or2b_1 _21355_ (.A(_14459_),
    .B_N(_14464_),
    .X(_01556_));
 sky130_fd_sc_hd__nand2_1 _21356_ (.A(_14458_),
    .B(_14465_),
    .Y(_01557_));
 sky130_fd_sc_hd__buf_2 _21357_ (.A(_12413_),
    .X(_01558_));
 sky130_fd_sc_hd__a31o_2 _21358_ (.A1(_11447_),
    .A2(_01558_),
    .A3(_14463_),
    .B1(_14461_),
    .X(_01559_));
 sky130_fd_sc_hd__o21ba_1 _21359_ (.A1(_14477_),
    .A2(_14479_),
    .B1_N(_14478_),
    .X(_01560_));
 sky130_fd_sc_hd__a22oi_1 _21360_ (.A1(_11666_),
    .A2(_12278_),
    .B1(_13667_),
    .B2(_11557_),
    .Y(_01561_));
 sky130_fd_sc_hd__and4_1 _21361_ (.A(_11664_),
    .B(_11782_),
    .C(_13674_),
    .D(_12413_),
    .X(_01562_));
 sky130_fd_sc_hd__nor2_1 _21362_ (.A(_01561_),
    .B(_01562_),
    .Y(_01563_));
 sky130_fd_sc_hd__clkbuf_2 _21363_ (.A(_12543_),
    .X(_01564_));
 sky130_fd_sc_hd__nand2_1 _21364_ (.A(_11561_),
    .B(_01564_),
    .Y(_01565_));
 sky130_fd_sc_hd__xnor2_2 _21365_ (.A(_01563_),
    .B(_01565_),
    .Y(_01566_));
 sky130_fd_sc_hd__xnor2_1 _21366_ (.A(_01560_),
    .B(_01566_),
    .Y(_01567_));
 sky130_fd_sc_hd__xnor2_1 _21367_ (.A(_01559_),
    .B(_01567_),
    .Y(_01568_));
 sky130_fd_sc_hd__a21oi_1 _21368_ (.A1(_01556_),
    .A2(_01557_),
    .B1(_01568_),
    .Y(_01569_));
 sky130_fd_sc_hd__and3_1 _21369_ (.A(_01556_),
    .B(_01557_),
    .C(_01568_),
    .X(_01570_));
 sky130_fd_sc_hd__nor3_1 _21370_ (.A(_01555_),
    .B(_01569_),
    .C(_01570_),
    .Y(_01571_));
 sky130_fd_sc_hd__o21a_1 _21371_ (.A1(_01569_),
    .A2(_01570_),
    .B1(_01555_),
    .X(_01572_));
 sky130_fd_sc_hd__a211o_1 _21372_ (.A1(_01536_),
    .A2(_14493_),
    .B1(net356),
    .C1(_01572_),
    .X(_01573_));
 sky130_fd_sc_hd__o211ai_1 _21373_ (.A1(net356),
    .A2(_01572_),
    .B1(_01536_),
    .C1(_14493_),
    .Y(_01574_));
 sky130_fd_sc_hd__nand2_1 _21374_ (.A(_01573_),
    .B(_01574_),
    .Y(_01575_));
 sky130_fd_sc_hd__xor2_1 _21375_ (.A(_01535_),
    .B(_01575_),
    .X(_01576_));
 sky130_fd_sc_hd__or2b_1 _21376_ (.A(_14488_),
    .B_N(_14487_),
    .X(_01577_));
 sky130_fd_sc_hd__nand2_1 _21377_ (.A(_14481_),
    .B(_14489_),
    .Y(_01578_));
 sky130_fd_sc_hd__or3_2 _21378_ (.A(_14496_),
    .B(_14500_),
    .C(_14501_),
    .X(_01579_));
 sky130_fd_sc_hd__nand2_1 _21379_ (.A(_11772_),
    .B(_14283_),
    .Y(_01580_));
 sky130_fd_sc_hd__and4_1 _21380_ (.A(_11954_),
    .B(_12075_),
    .C(_13936_),
    .D(_13937_),
    .X(_01581_));
 sky130_fd_sc_hd__buf_2 _21381_ (.A(_13713_),
    .X(_01582_));
 sky130_fd_sc_hd__buf_4 _21382_ (.A(_13716_),
    .X(_01583_));
 sky130_fd_sc_hd__a22oi_1 _21383_ (.A1(_13919_),
    .A2(_01582_),
    .B1(_01583_),
    .B2(_11954_),
    .Y(_01584_));
 sky130_fd_sc_hd__nor2_1 _21384_ (.A(_01581_),
    .B(_01584_),
    .Y(_01585_));
 sky130_fd_sc_hd__xnor2_2 _21385_ (.A(_01580_),
    .B(_01585_),
    .Y(_01586_));
 sky130_fd_sc_hd__nand2_1 _21386_ (.A(_11826_),
    .B(_13720_),
    .Y(_01587_));
 sky130_fd_sc_hd__and4_1 _21387_ (.A(_12343_),
    .B(_12561_),
    .C(_12329_),
    .D(_14129_),
    .X(_01588_));
 sky130_fd_sc_hd__a22oi_2 _21388_ (.A1(_11381_),
    .A2(_14132_),
    .B1(_14310_),
    .B2(_11373_),
    .Y(_01589_));
 sky130_fd_sc_hd__nor2_1 _21389_ (.A(_01588_),
    .B(_01589_),
    .Y(_01590_));
 sky130_fd_sc_hd__xnor2_1 _21390_ (.A(_01587_),
    .B(_01590_),
    .Y(_01591_));
 sky130_fd_sc_hd__o21ba_1 _21391_ (.A1(_14483_),
    .A2(_14485_),
    .B1_N(_14484_),
    .X(_01592_));
 sky130_fd_sc_hd__xnor2_1 _21392_ (.A(_01591_),
    .B(_01592_),
    .Y(_01593_));
 sky130_fd_sc_hd__xnor2_1 _21393_ (.A(_01586_),
    .B(_01593_),
    .Y(_01594_));
 sky130_fd_sc_hd__a21oi_1 _21394_ (.A1(_01579_),
    .A2(_14504_),
    .B1(_01594_),
    .Y(_01595_));
 sky130_fd_sc_hd__and3_1 _21395_ (.A(_01579_),
    .B(_14504_),
    .C(_01594_),
    .X(_01596_));
 sky130_fd_sc_hd__a211o_1 _21396_ (.A1(_01577_),
    .A2(_01578_),
    .B1(_01595_),
    .C1(_01596_),
    .X(_01597_));
 sky130_fd_sc_hd__o211ai_1 _21397_ (.A1(_01595_),
    .A2(_01596_),
    .B1(_01577_),
    .C1(_01578_),
    .Y(_01598_));
 sky130_fd_sc_hd__and2_1 _21398_ (.A(_01597_),
    .B(_01598_),
    .X(_01599_));
 sky130_fd_sc_hd__o21ba_1 _21399_ (.A1(_14507_),
    .A2(_14511_),
    .B1_N(_14509_),
    .X(_01600_));
 sky130_fd_sc_hd__buf_2 _21400_ (.A(_12910_),
    .X(_01601_));
 sky130_fd_sc_hd__and4_2 _21401_ (.A(_11269_),
    .B(_11055_),
    .C(_12771_),
    .D(_01601_),
    .X(_01602_));
 sky130_fd_sc_hd__a22oi_1 _21402_ (.A1(_11728_),
    .A2(_13743_),
    .B1(_13741_),
    .B2(_11043_),
    .Y(_01603_));
 sky130_fd_sc_hd__and4bb_1 _21403_ (.A_N(_01602_),
    .B_N(_01603_),
    .C(_11262_),
    .D(_14147_),
    .X(_01604_));
 sky130_fd_sc_hd__o2bb2a_1 _21404_ (.A1_N(_11474_),
    .A2_N(_13738_),
    .B1(_01602_),
    .B2(_01603_),
    .X(_01605_));
 sky130_fd_sc_hd__nor2_1 _21405_ (.A(_01604_),
    .B(_01605_),
    .Y(_01606_));
 sky130_fd_sc_hd__xnor2_1 _21406_ (.A(_01600_),
    .B(_01606_),
    .Y(_01607_));
 sky130_fd_sc_hd__o21ai_2 _21407_ (.A1(_14497_),
    .A2(_14500_),
    .B1(_01607_),
    .Y(_01608_));
 sky130_fd_sc_hd__or3_1 _21408_ (.A(_14497_),
    .B(_14500_),
    .C(_01607_),
    .X(_01609_));
 sky130_fd_sc_hd__and2_1 _21409_ (.A(_01608_),
    .B(_01609_),
    .X(_01610_));
 sky130_fd_sc_hd__nand2_1 _21410_ (.A(_11167_),
    .B(_13226_),
    .Y(_01611_));
 sky130_fd_sc_hd__and4_1 _21411_ (.A(_11405_),
    .B(_11402_),
    .C(_13761_),
    .D(_13762_),
    .X(_01612_));
 sky130_fd_sc_hd__clkbuf_4 _21412_ (.A(_13765_),
    .X(_01613_));
 sky130_fd_sc_hd__a22oi_2 _21413_ (.A1(_11402_),
    .A2(_13224_),
    .B1(_01613_),
    .B2(_13959_),
    .Y(_01614_));
 sky130_fd_sc_hd__nor2_1 _21414_ (.A(_01612_),
    .B(_01614_),
    .Y(_01615_));
 sky130_fd_sc_hd__xnor2_2 _21415_ (.A(_01611_),
    .B(_01615_),
    .Y(_01616_));
 sky130_fd_sc_hd__nand2_1 _21416_ (.A(_12361_),
    .B(_13752_),
    .Y(_01617_));
 sky130_fd_sc_hd__buf_2 _21417_ (.A(\genblk1.pcpi_mul.rs2[32] ),
    .X(_01618_));
 sky130_fd_sc_hd__and2b_1 _21418_ (.A_N(_10742_),
    .B(_01618_),
    .X(_01619_));
 sky130_fd_sc_hd__clkbuf_2 _21419_ (.A(\genblk1.pcpi_mul.rs2[31] ),
    .X(_01620_));
 sky130_fd_sc_hd__nand2_1 _21420_ (.A(_11199_),
    .B(_01620_),
    .Y(_01621_));
 sky130_fd_sc_hd__xnor2_2 _21421_ (.A(_01619_),
    .B(_01621_),
    .Y(_01622_));
 sky130_fd_sc_hd__xnor2_2 _21422_ (.A(_01617_),
    .B(_01622_),
    .Y(_01623_));
 sky130_fd_sc_hd__buf_2 _21423_ (.A(_14342_),
    .X(_01624_));
 sky130_fd_sc_hd__buf_2 _21424_ (.A(_13753_),
    .X(_01625_));
 sky130_fd_sc_hd__and3_1 _21425_ (.A(_11245_),
    .B(_01625_),
    .C(_14515_),
    .X(_01626_));
 sky130_fd_sc_hd__a31o_2 _21426_ (.A1(_11343_),
    .A2(_01624_),
    .A3(_14517_),
    .B1(_01626_),
    .X(_01627_));
 sky130_fd_sc_hd__xor2_2 _21427_ (.A(_01623_),
    .B(_01627_),
    .X(_01628_));
 sky130_fd_sc_hd__xnor2_1 _21428_ (.A(_01616_),
    .B(_01628_),
    .Y(_01629_));
 sky130_fd_sc_hd__nand2_1 _21429_ (.A(_14518_),
    .B(_14520_),
    .Y(_01630_));
 sky130_fd_sc_hd__a21boi_2 _21430_ (.A1(_14513_),
    .A2(_14521_),
    .B1_N(_01630_),
    .Y(_01631_));
 sky130_fd_sc_hd__xnor2_1 _21431_ (.A(_01629_),
    .B(_01631_),
    .Y(_01632_));
 sky130_fd_sc_hd__xnor2_1 _21432_ (.A(_01610_),
    .B(_01632_),
    .Y(_01633_));
 sky130_fd_sc_hd__nand2_1 _21433_ (.A(_14522_),
    .B(_14524_),
    .Y(_01634_));
 sky130_fd_sc_hd__nor2_1 _21434_ (.A(_14522_),
    .B(_14524_),
    .Y(_01635_));
 sky130_fd_sc_hd__a21oi_1 _21435_ (.A1(_14506_),
    .A2(_01634_),
    .B1(_01635_),
    .Y(_01636_));
 sky130_fd_sc_hd__xnor2_1 _21436_ (.A(_01633_),
    .B(_01636_),
    .Y(_01637_));
 sky130_fd_sc_hd__xnor2_1 _21437_ (.A(_01599_),
    .B(_01637_),
    .Y(_01638_));
 sky130_fd_sc_hd__and2b_1 _21438_ (.A_N(_14529_),
    .B(_14526_),
    .X(_01639_));
 sky130_fd_sc_hd__a21oi_2 _21439_ (.A1(_14495_),
    .A2(_14530_),
    .B1(_01639_),
    .Y(_01640_));
 sky130_fd_sc_hd__xor2_1 _21440_ (.A(_01638_),
    .B(_01640_),
    .X(_01641_));
 sky130_fd_sc_hd__xor2_1 _21441_ (.A(_01576_),
    .B(_01641_),
    .X(_01642_));
 sky130_fd_sc_hd__nor2_1 _21442_ (.A(_14531_),
    .B(_14533_),
    .Y(_01643_));
 sky130_fd_sc_hd__a21oi_2 _21443_ (.A1(_14473_),
    .A2(_14534_),
    .B1(_01643_),
    .Y(_01644_));
 sky130_fd_sc_hd__xnor2_1 _21444_ (.A(_01642_),
    .B(_01644_),
    .Y(_01645_));
 sky130_fd_sc_hd__xor2_1 _21445_ (.A(_01534_),
    .B(_01645_),
    .X(_01646_));
 sky130_fd_sc_hd__and2b_1 _21446_ (.A_N(_14537_),
    .B(_14535_),
    .X(_01647_));
 sky130_fd_sc_hd__a21oi_4 _21447_ (.A1(_14435_),
    .A2(_14538_),
    .B1(_01647_),
    .Y(_01648_));
 sky130_fd_sc_hd__xnor2_1 _21448_ (.A(_01646_),
    .B(_01648_),
    .Y(_01649_));
 sky130_fd_sc_hd__xnor2_1 _21449_ (.A(_14557_),
    .B(_01649_),
    .Y(_01650_));
 sky130_fd_sc_hd__nor2_1 _21450_ (.A(_14539_),
    .B(_14541_),
    .Y(_01651_));
 sky130_fd_sc_hd__a21oi_4 _21451_ (.A1(_14387_),
    .A2(_14542_),
    .B1(_01651_),
    .Y(_01652_));
 sky130_fd_sc_hd__xor2_1 _21452_ (.A(_01650_),
    .B(_01652_),
    .X(_01653_));
 sky130_fd_sc_hd__xnor2_1 _21453_ (.A(_14385_),
    .B(_01653_),
    .Y(_01654_));
 sky130_fd_sc_hd__nor2_1 _21454_ (.A(_14543_),
    .B(_14545_),
    .Y(_01655_));
 sky130_fd_sc_hd__a21oi_4 _21455_ (.A1(_14381_),
    .A2(_14546_),
    .B1(_01655_),
    .Y(_01656_));
 sky130_fd_sc_hd__or2_1 _21456_ (.A(_01654_),
    .B(_01656_),
    .X(_01657_));
 sky130_fd_sc_hd__nand2_1 _21457_ (.A(_01654_),
    .B(_01656_),
    .Y(_01658_));
 sky130_fd_sc_hd__nand2_2 _21458_ (.A(_01657_),
    .B(_01658_),
    .Y(_01659_));
 sky130_fd_sc_hd__nand2_1 _21459_ (.A(_14380_),
    .B(_14547_),
    .Y(_01660_));
 sky130_fd_sc_hd__and2b_2 _21460_ (.A_N(_14375_),
    .B(_14548_),
    .X(_01661_));
 sky130_fd_sc_hd__nor2_1 _21461_ (.A(_14380_),
    .B(_14547_),
    .Y(_01662_));
 sky130_fd_sc_hd__a221oi_4 _21462_ (.A1(_14550_),
    .A2(_01660_),
    .B1(_01661_),
    .B2(_14377_),
    .C1(_01662_),
    .Y(_01663_));
 sky130_fd_sc_hd__nand2_4 _21463_ (.A(_14376_),
    .B(_01661_),
    .Y(_01664_));
 sky130_fd_sc_hd__a21o_1 _21464_ (.A1(_14007_),
    .A2(_14009_),
    .B1(_01664_),
    .X(_01665_));
 sky130_fd_sc_hd__nand2_2 _21465_ (.A(net334),
    .B(_01665_),
    .Y(_01666_));
 sky130_fd_sc_hd__xnor2_4 _21466_ (.A(_01659_),
    .B(_01666_),
    .Y(_00082_));
 sky130_fd_sc_hd__nor2_1 _21467_ (.A(_01650_),
    .B(_01652_),
    .Y(_01667_));
 sky130_fd_sc_hd__a21o_1 _21468_ (.A1(_14385_),
    .A2(_01653_),
    .B1(_01667_),
    .X(_01668_));
 sky130_fd_sc_hd__and2b_1 _21469_ (.A_N(_01532_),
    .B(_14561_),
    .X(_01669_));
 sky130_fd_sc_hd__and2b_1 _21470_ (.A_N(_14559_),
    .B(_01533_),
    .X(_01670_));
 sky130_fd_sc_hd__a21oi_1 _21471_ (.A1(_14567_),
    .A2(_01509_),
    .B1(_01507_),
    .Y(_01671_));
 sky130_fd_sc_hd__o21ba_2 _21472_ (.A1(_01669_),
    .A2(_01670_),
    .B1_N(_01671_),
    .X(_01672_));
 sky130_fd_sc_hd__or3b_1 _21473_ (.A(_01669_),
    .B(_01670_),
    .C_N(_01671_),
    .X(_01673_));
 sky130_fd_sc_hd__and2b_1 _21474_ (.A_N(_01672_),
    .B(_01673_),
    .X(_01674_));
 sky130_fd_sc_hd__o32a_1 _21475_ (.A1(_01526_),
    .A2(_01527_),
    .A3(_01530_),
    .B1(_01531_),
    .B2(_01510_),
    .X(_01675_));
 sky130_fd_sc_hd__o21a_1 _21476_ (.A1(_01535_),
    .A2(_01575_),
    .B1(_01573_),
    .X(_01676_));
 sky130_fd_sc_hd__nand2_1 _21477_ (.A(_14569_),
    .B(_01502_),
    .Y(_01677_));
 sky130_fd_sc_hd__and3_1 _21478_ (.A(_10663_),
    .B(_14223_),
    .C(_14038_),
    .X(_01678_));
 sky130_fd_sc_hd__o21ai_4 _21479_ (.A1(_10663_),
    .A2(_14223_),
    .B1(_14563_),
    .Y(_01679_));
 sky130_fd_sc_hd__nor2_1 _21480_ (.A(_01678_),
    .B(_01679_),
    .Y(_01680_));
 sky130_fd_sc_hd__o22a_2 _21481_ (.A1(_14222_),
    .A2(_14571_),
    .B1(_01500_),
    .B2(_10585_),
    .X(_01681_));
 sky130_fd_sc_hd__xnor2_2 _21482_ (.A(_01680_),
    .B(_01681_),
    .Y(_01682_));
 sky130_fd_sc_hd__xor2_1 _21483_ (.A(_14395_),
    .B(_01682_),
    .X(_01683_));
 sky130_fd_sc_hd__a21oi_2 _21484_ (.A1(_01677_),
    .A2(_01504_),
    .B1(_01683_),
    .Y(_01684_));
 sky130_fd_sc_hd__and3_1 _21485_ (.A(_01677_),
    .B(_01504_),
    .C(_01683_),
    .X(_01685_));
 sky130_fd_sc_hd__nor2_1 _21486_ (.A(_01684_),
    .B(_01685_),
    .Y(_01686_));
 sky130_fd_sc_hd__xnor2_1 _21487_ (.A(_14567_),
    .B(_01686_),
    .Y(_01687_));
 sky130_fd_sc_hd__or2b_1 _21488_ (.A(_01515_),
    .B_N(_01521_),
    .X(_01688_));
 sky130_fd_sc_hd__or2b_1 _21489_ (.A(_01514_),
    .B_N(_01522_),
    .X(_01689_));
 sky130_fd_sc_hd__nand2_1 _21490_ (.A(_01688_),
    .B(_01689_),
    .Y(_01690_));
 sky130_fd_sc_hd__and2b_1 _21491_ (.A_N(_01551_),
    .B(_01550_),
    .X(_01691_));
 sky130_fd_sc_hd__o21ba_1 _21492_ (.A1(_01517_),
    .A2(_01520_),
    .B1_N(_01518_),
    .X(_01692_));
 sky130_fd_sc_hd__o21ba_1 _21493_ (.A1(_01537_),
    .A2(_01541_),
    .B1_N(_01539_),
    .X(_01693_));
 sky130_fd_sc_hd__a22oi_1 _21494_ (.A1(_13858_),
    .A2(_13824_),
    .B1(_13826_),
    .B2(_10784_),
    .Y(_01694_));
 sky130_fd_sc_hd__and4_1 _21495_ (.A(_13863_),
    .B(_14055_),
    .C(_14033_),
    .D(_13606_),
    .X(_01695_));
 sky130_fd_sc_hd__nor2_1 _21496_ (.A(_01694_),
    .B(_01695_),
    .Y(_01696_));
 sky130_fd_sc_hd__nand2_1 _21497_ (.A(_10738_),
    .B(_14211_),
    .Y(_01697_));
 sky130_fd_sc_hd__xnor2_1 _21498_ (.A(_01696_),
    .B(_01697_),
    .Y(_01698_));
 sky130_fd_sc_hd__xnor2_1 _21499_ (.A(_01693_),
    .B(_01698_),
    .Y(_01699_));
 sky130_fd_sc_hd__xnor2_2 _21500_ (.A(_01692_),
    .B(_01699_),
    .Y(_01700_));
 sky130_fd_sc_hd__o21ai_2 _21501_ (.A1(_01691_),
    .A2(_01553_),
    .B1(_01700_),
    .Y(_01701_));
 sky130_fd_sc_hd__or3_1 _21502_ (.A(_01691_),
    .B(_01553_),
    .C(_01700_),
    .X(_01702_));
 sky130_fd_sc_hd__nand3_1 _21503_ (.A(_01690_),
    .B(_01701_),
    .C(_01702_),
    .Y(_01703_));
 sky130_fd_sc_hd__a21o_1 _21504_ (.A1(_01701_),
    .A2(_01702_),
    .B1(_01690_),
    .X(_01704_));
 sky130_fd_sc_hd__o211a_1 _21505_ (.A1(_01524_),
    .A2(_01526_),
    .B1(_01703_),
    .C1(_01704_),
    .X(_01705_));
 sky130_fd_sc_hd__a211oi_1 _21506_ (.A1(_01703_),
    .A2(_01704_),
    .B1(_01524_),
    .C1(_01526_),
    .Y(_01706_));
 sky130_fd_sc_hd__nor2_1 _21507_ (.A(_01705_),
    .B(_01706_),
    .Y(_01707_));
 sky130_fd_sc_hd__xnor2_1 _21508_ (.A(_01687_),
    .B(_01707_),
    .Y(_01708_));
 sky130_fd_sc_hd__xnor2_1 _21509_ (.A(_01676_),
    .B(_01708_),
    .Y(_01709_));
 sky130_fd_sc_hd__xnor2_2 _21510_ (.A(_01675_),
    .B(_01709_),
    .Y(_01710_));
 sky130_fd_sc_hd__nor2_2 _21511_ (.A(_01569_),
    .B(_01571_),
    .Y(_01711_));
 sky130_fd_sc_hd__a21o_1 _21512_ (.A1(_01579_),
    .A2(_14504_),
    .B1(_01594_),
    .X(_01712_));
 sky130_fd_sc_hd__clkbuf_2 _21513_ (.A(_13445_),
    .X(_01713_));
 sky130_fd_sc_hd__a22oi_1 _21514_ (.A1(_13662_),
    .A2(_13868_),
    .B1(_01713_),
    .B2(_13661_),
    .Y(_01714_));
 sky130_fd_sc_hd__and4_1 _21515_ (.A(_13669_),
    .B(_11112_),
    .C(_13285_),
    .D(_14417_),
    .X(_01715_));
 sky130_fd_sc_hd__nor2_1 _21516_ (.A(_01714_),
    .B(_01715_),
    .Y(_01716_));
 sky130_fd_sc_hd__buf_2 _21517_ (.A(_01516_),
    .X(_01717_));
 sky130_fd_sc_hd__clkbuf_2 _21518_ (.A(_01717_),
    .X(_01718_));
 sky130_fd_sc_hd__nand2_1 _21519_ (.A(_10895_),
    .B(_01718_),
    .Y(_01719_));
 sky130_fd_sc_hd__xnor2_2 _21520_ (.A(_01716_),
    .B(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__nand2_1 _21521_ (.A(_11233_),
    .B(_14262_),
    .Y(_01721_));
 sky130_fd_sc_hd__and4_1 _21522_ (.A(_13899_),
    .B(_13900_),
    .C(_14080_),
    .D(_14076_),
    .X(_01722_));
 sky130_fd_sc_hd__a22oi_2 _21523_ (.A1(_13903_),
    .A2(_14444_),
    .B1(_13860_),
    .B2(_11242_),
    .Y(_01723_));
 sky130_fd_sc_hd__nor2_1 _21524_ (.A(_01722_),
    .B(_01723_),
    .Y(_01724_));
 sky130_fd_sc_hd__xnor2_2 _21525_ (.A(_01721_),
    .B(_01724_),
    .Y(_01725_));
 sky130_fd_sc_hd__o21ba_1 _21526_ (.A1(_01545_),
    .A2(_01548_),
    .B1_N(_01546_),
    .X(_01726_));
 sky130_fd_sc_hd__xnor2_1 _21527_ (.A(_01725_),
    .B(_01726_),
    .Y(_01727_));
 sky130_fd_sc_hd__and2_1 _21528_ (.A(_01720_),
    .B(_01727_),
    .X(_01728_));
 sky130_fd_sc_hd__nor2_1 _21529_ (.A(_01720_),
    .B(_01727_),
    .Y(_01729_));
 sky130_fd_sc_hd__or2_2 _21530_ (.A(_01728_),
    .B(_01729_),
    .X(_01730_));
 sky130_fd_sc_hd__or2b_1 _21531_ (.A(_01560_),
    .B_N(_01566_),
    .X(_01731_));
 sky130_fd_sc_hd__nand2_1 _21532_ (.A(_01559_),
    .B(_01567_),
    .Y(_01732_));
 sky130_fd_sc_hd__a31o_2 _21533_ (.A1(_11447_),
    .A2(_01564_),
    .A3(_01563_),
    .B1(_01562_),
    .X(_01733_));
 sky130_fd_sc_hd__o21ba_2 _21534_ (.A1(_01580_),
    .A2(_01584_),
    .B1_N(_01581_),
    .X(_01734_));
 sky130_fd_sc_hd__a22oi_1 _21535_ (.A1(_11666_),
    .A2(_12413_),
    .B1(_13668_),
    .B2(_11557_),
    .Y(_01735_));
 sky130_fd_sc_hd__and4_1 _21536_ (.A(_14105_),
    .B(_11782_),
    .C(_13666_),
    .D(_13484_),
    .X(_01736_));
 sky130_fd_sc_hd__nor2_1 _21537_ (.A(_01735_),
    .B(_01736_),
    .Y(_01737_));
 sky130_fd_sc_hd__nand2_1 _21538_ (.A(_11561_),
    .B(_13659_),
    .Y(_01738_));
 sky130_fd_sc_hd__xnor2_2 _21539_ (.A(_01737_),
    .B(_01738_),
    .Y(_01739_));
 sky130_fd_sc_hd__xnor2_1 _21540_ (.A(_01734_),
    .B(_01739_),
    .Y(_01740_));
 sky130_fd_sc_hd__xnor2_1 _21541_ (.A(_01733_),
    .B(_01740_),
    .Y(_01741_));
 sky130_fd_sc_hd__a21oi_1 _21542_ (.A1(_01731_),
    .A2(_01732_),
    .B1(_01741_),
    .Y(_01742_));
 sky130_fd_sc_hd__and3_1 _21543_ (.A(_01731_),
    .B(_01732_),
    .C(_01741_),
    .X(_01743_));
 sky130_fd_sc_hd__nor3_1 _21544_ (.A(_01730_),
    .B(_01742_),
    .C(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__o21a_1 _21545_ (.A1(_01742_),
    .A2(_01743_),
    .B1(_01730_),
    .X(_01745_));
 sky130_fd_sc_hd__a211o_1 _21546_ (.A1(_01712_),
    .A2(_01597_),
    .B1(_01744_),
    .C1(_01745_),
    .X(_01746_));
 sky130_fd_sc_hd__o211ai_1 _21547_ (.A1(_01744_),
    .A2(_01745_),
    .B1(_01712_),
    .C1(_01597_),
    .Y(_01747_));
 sky130_fd_sc_hd__nand2_2 _21548_ (.A(_01746_),
    .B(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__xor2_2 _21549_ (.A(_01711_),
    .B(_01748_),
    .X(_01749_));
 sky130_fd_sc_hd__or2b_1 _21550_ (.A(_01592_),
    .B_N(_01591_),
    .X(_01750_));
 sky130_fd_sc_hd__nand2_1 _21551_ (.A(_01586_),
    .B(_01593_),
    .Y(_01751_));
 sky130_fd_sc_hd__or3_1 _21552_ (.A(_01600_),
    .B(_01604_),
    .C(_01605_),
    .X(_01752_));
 sky130_fd_sc_hd__nand2_1 _21553_ (.A(_13711_),
    .B(_14457_),
    .Y(_01753_));
 sky130_fd_sc_hd__buf_2 _21554_ (.A(_13713_),
    .X(_01754_));
 sky130_fd_sc_hd__buf_2 _21555_ (.A(_13715_),
    .X(_01755_));
 sky130_fd_sc_hd__and4_1 _21556_ (.A(_11820_),
    .B(_13904_),
    .C(_01754_),
    .D(_01755_),
    .X(_01756_));
 sky130_fd_sc_hd__buf_2 _21557_ (.A(_13715_),
    .X(_01757_));
 sky130_fd_sc_hd__a22oi_2 _21558_ (.A1(_13904_),
    .A2(_01582_),
    .B1(_01757_),
    .B2(_12075_),
    .Y(_01758_));
 sky130_fd_sc_hd__nor2_1 _21559_ (.A(_01756_),
    .B(_01758_),
    .Y(_01759_));
 sky130_fd_sc_hd__xnor2_2 _21560_ (.A(_01753_),
    .B(_01759_),
    .Y(_01760_));
 sky130_fd_sc_hd__nand2_1 _21561_ (.A(_13690_),
    .B(_12227_),
    .Y(_01761_));
 sky130_fd_sc_hd__and4_1 _21562_ (.A(_12561_),
    .B(_11490_),
    .C(_12323_),
    .D(_14129_),
    .X(_01762_));
 sky130_fd_sc_hd__a22oi_2 _21563_ (.A1(_11591_),
    .A2(_13942_),
    .B1(_14310_),
    .B2(_11381_),
    .Y(_01763_));
 sky130_fd_sc_hd__nor2_1 _21564_ (.A(_01762_),
    .B(_01763_),
    .Y(_01764_));
 sky130_fd_sc_hd__xnor2_1 _21565_ (.A(_01761_),
    .B(_01764_),
    .Y(_01765_));
 sky130_fd_sc_hd__o21ba_1 _21566_ (.A1(_01587_),
    .A2(_01589_),
    .B1_N(_01588_),
    .X(_01766_));
 sky130_fd_sc_hd__xnor2_1 _21567_ (.A(_01765_),
    .B(_01766_),
    .Y(_01767_));
 sky130_fd_sc_hd__xnor2_1 _21568_ (.A(_01760_),
    .B(_01767_),
    .Y(_01768_));
 sky130_fd_sc_hd__a21oi_1 _21569_ (.A1(_01752_),
    .A2(_01608_),
    .B1(_01768_),
    .Y(_01769_));
 sky130_fd_sc_hd__and3_1 _21570_ (.A(_01752_),
    .B(_01608_),
    .C(_01768_),
    .X(_01770_));
 sky130_fd_sc_hd__a211o_1 _21571_ (.A1(_01750_),
    .A2(_01751_),
    .B1(_01769_),
    .C1(_01770_),
    .X(_01771_));
 sky130_fd_sc_hd__o211ai_1 _21572_ (.A1(_01769_),
    .A2(_01770_),
    .B1(_01750_),
    .C1(_01751_),
    .Y(_01772_));
 sky130_fd_sc_hd__and2_1 _21573_ (.A(_01771_),
    .B(_01772_),
    .X(_01773_));
 sky130_fd_sc_hd__o21ba_1 _21574_ (.A1(_01611_),
    .A2(_01614_),
    .B1_N(_01612_),
    .X(_01774_));
 sky130_fd_sc_hd__and4_1 _21575_ (.A(_11055_),
    .B(_11601_),
    .C(_12776_),
    .D(_01601_),
    .X(_01775_));
 sky130_fd_sc_hd__a22oi_1 _21576_ (.A1(_11473_),
    .A2(_13743_),
    .B1(_13741_),
    .B2(_11728_),
    .Y(_01776_));
 sky130_fd_sc_hd__and4bb_1 _21577_ (.A_N(_01775_),
    .B_N(_01776_),
    .C(_11278_),
    .D(_14147_),
    .X(_01777_));
 sky130_fd_sc_hd__o2bb2a_1 _21578_ (.A1_N(_11369_),
    .A2_N(_13738_),
    .B1(_01775_),
    .B2(_01776_),
    .X(_01778_));
 sky130_fd_sc_hd__nor2_1 _21579_ (.A(_01777_),
    .B(_01778_),
    .Y(_01779_));
 sky130_fd_sc_hd__xnor2_1 _21580_ (.A(_01774_),
    .B(_01779_),
    .Y(_01780_));
 sky130_fd_sc_hd__o21ai_2 _21581_ (.A1(_01602_),
    .A2(_01604_),
    .B1(_01780_),
    .Y(_01781_));
 sky130_fd_sc_hd__or3_1 _21582_ (.A(_01602_),
    .B(_01604_),
    .C(_01780_),
    .X(_01782_));
 sky130_fd_sc_hd__and2_1 _21583_ (.A(_01781_),
    .B(_01782_),
    .X(_01783_));
 sky130_fd_sc_hd__nand2_1 _21584_ (.A(_11157_),
    .B(_13226_),
    .Y(_01784_));
 sky130_fd_sc_hd__and4_1 _21585_ (.A(_11049_),
    .B(_11037_),
    .C(_13761_),
    .D(_14508_),
    .X(_01785_));
 sky130_fd_sc_hd__a22oi_2 _21586_ (.A1(_11386_),
    .A2(_13970_),
    .B1(_14510_),
    .B2(_11402_),
    .Y(_01786_));
 sky130_fd_sc_hd__nor2_1 _21587_ (.A(_01785_),
    .B(_01786_),
    .Y(_01787_));
 sky130_fd_sc_hd__xnor2_2 _21588_ (.A(_01784_),
    .B(_01787_),
    .Y(_01788_));
 sky130_fd_sc_hd__nand2_1 _21589_ (.A(_13959_),
    .B(_13752_),
    .Y(_01789_));
 sky130_fd_sc_hd__and2b_1 _21590_ (.A_N(_10746_),
    .B(_01618_),
    .X(_01790_));
 sky130_fd_sc_hd__nand2_1 _21591_ (.A(_11302_),
    .B(_13753_),
    .Y(_01791_));
 sky130_fd_sc_hd__xnor2_2 _21592_ (.A(_01790_),
    .B(_01791_),
    .Y(_01792_));
 sky130_fd_sc_hd__xnor2_2 _21593_ (.A(_01789_),
    .B(_01792_),
    .Y(_01793_));
 sky130_fd_sc_hd__and3_1 _21594_ (.A(_11343_),
    .B(_01625_),
    .C(_01619_),
    .X(_01794_));
 sky130_fd_sc_hd__a31o_2 _21595_ (.A1(_12361_),
    .A2(_01624_),
    .A3(_01622_),
    .B1(_01794_),
    .X(_01795_));
 sky130_fd_sc_hd__xor2_2 _21596_ (.A(_01793_),
    .B(_01795_),
    .X(_01796_));
 sky130_fd_sc_hd__xnor2_2 _21597_ (.A(_01788_),
    .B(_01796_),
    .Y(_01797_));
 sky130_fd_sc_hd__nand2_1 _21598_ (.A(_01623_),
    .B(_01627_),
    .Y(_01798_));
 sky130_fd_sc_hd__a21boi_2 _21599_ (.A1(_01616_),
    .A2(_01628_),
    .B1_N(_01798_),
    .Y(_01799_));
 sky130_fd_sc_hd__xnor2_1 _21600_ (.A(_01797_),
    .B(_01799_),
    .Y(_01800_));
 sky130_fd_sc_hd__xnor2_2 _21601_ (.A(_01783_),
    .B(_01800_),
    .Y(_01801_));
 sky130_fd_sc_hd__nand2_1 _21602_ (.A(_01629_),
    .B(_01631_),
    .Y(_01802_));
 sky130_fd_sc_hd__nor2_1 _21603_ (.A(_01629_),
    .B(_01631_),
    .Y(_01803_));
 sky130_fd_sc_hd__a21oi_2 _21604_ (.A1(_01610_),
    .A2(_01802_),
    .B1(_01803_),
    .Y(_01804_));
 sky130_fd_sc_hd__xnor2_2 _21605_ (.A(_01801_),
    .B(_01804_),
    .Y(_01805_));
 sky130_fd_sc_hd__xnor2_2 _21606_ (.A(_01773_),
    .B(_01805_),
    .Y(_01806_));
 sky130_fd_sc_hd__and2b_1 _21607_ (.A_N(_01636_),
    .B(_01633_),
    .X(_01807_));
 sky130_fd_sc_hd__a21oi_2 _21608_ (.A1(_01599_),
    .A2(_01637_),
    .B1(_01807_),
    .Y(_01808_));
 sky130_fd_sc_hd__xor2_2 _21609_ (.A(_01806_),
    .B(_01808_),
    .X(_01809_));
 sky130_fd_sc_hd__xor2_2 _21610_ (.A(_01749_),
    .B(_01809_),
    .X(_01810_));
 sky130_fd_sc_hd__nor2_1 _21611_ (.A(_01638_),
    .B(_01640_),
    .Y(_01811_));
 sky130_fd_sc_hd__a21oi_2 _21612_ (.A1(_01576_),
    .A2(_01641_),
    .B1(_01811_),
    .Y(_01812_));
 sky130_fd_sc_hd__xnor2_2 _21613_ (.A(_01810_),
    .B(_01812_),
    .Y(_01813_));
 sky130_fd_sc_hd__xor2_2 _21614_ (.A(_01710_),
    .B(_01813_),
    .X(_01814_));
 sky130_fd_sc_hd__and2b_1 _21615_ (.A_N(_01644_),
    .B(_01642_),
    .X(_01815_));
 sky130_fd_sc_hd__a21oi_2 _21616_ (.A1(_01534_),
    .A2(_01645_),
    .B1(_01815_),
    .Y(_01816_));
 sky130_fd_sc_hd__xnor2_2 _21617_ (.A(_01814_),
    .B(_01816_),
    .Y(_01817_));
 sky130_fd_sc_hd__xnor2_1 _21618_ (.A(_01674_),
    .B(_01817_),
    .Y(_01818_));
 sky130_fd_sc_hd__or2b_1 _21619_ (.A(_01648_),
    .B_N(_01646_),
    .X(_01819_));
 sky130_fd_sc_hd__a21boi_1 _21620_ (.A1(_14557_),
    .A2(_01649_),
    .B1_N(_01819_),
    .Y(_01820_));
 sky130_fd_sc_hd__xor2_1 _21621_ (.A(_01818_),
    .B(_01820_),
    .X(_01821_));
 sky130_fd_sc_hd__xor2_1 _21622_ (.A(_14555_),
    .B(_01821_),
    .X(_01822_));
 sky130_fd_sc_hd__nand2_1 _21623_ (.A(_01668_),
    .B(_01822_),
    .Y(_01823_));
 sky130_fd_sc_hd__or2_1 _21624_ (.A(_01668_),
    .B(_01822_),
    .X(_01824_));
 sky130_fd_sc_hd__and2_2 _21625_ (.A(_01823_),
    .B(_01824_),
    .X(_01825_));
 sky130_fd_sc_hd__a21bo_1 _21626_ (.A1(_01658_),
    .A2(_01666_),
    .B1_N(_01657_),
    .X(_01826_));
 sky130_fd_sc_hd__xor2_4 _21627_ (.A(_01825_),
    .B(_01826_),
    .X(_00083_));
 sky130_fd_sc_hd__and2b_1 _21628_ (.A_N(_01676_),
    .B(_01708_),
    .X(_01827_));
 sky130_fd_sc_hd__and2b_1 _21629_ (.A_N(_01675_),
    .B(_01709_),
    .X(_01828_));
 sky130_fd_sc_hd__nor2_2 _21630_ (.A(_01827_),
    .B(_01828_),
    .Y(_01829_));
 sky130_fd_sc_hd__a21oi_4 _21631_ (.A1(_14567_),
    .A2(_01686_),
    .B1(_01684_),
    .Y(_01830_));
 sky130_fd_sc_hd__xnor2_4 _21632_ (.A(_01829_),
    .B(_01830_),
    .Y(_01831_));
 sky130_fd_sc_hd__o21ba_1 _21633_ (.A1(_01687_),
    .A2(_01706_),
    .B1_N(_01705_),
    .X(_01832_));
 sky130_fd_sc_hd__o21ai_4 _21634_ (.A1(_01711_),
    .A2(_01748_),
    .B1(_01746_),
    .Y(_01833_));
 sky130_fd_sc_hd__nand2_1 _21635_ (.A(_14222_),
    .B(_01679_),
    .Y(_01834_));
 sky130_fd_sc_hd__xnor2_1 _21636_ (.A(_14395_),
    .B(_01834_),
    .Y(_01835_));
 sky130_fd_sc_hd__o21a_1 _21637_ (.A1(_01682_),
    .A2(_01835_),
    .B1(_14566_),
    .X(_01836_));
 sky130_fd_sc_hd__nor3_1 _21638_ (.A(_14567_),
    .B(_01682_),
    .C(_01835_),
    .Y(_01837_));
 sky130_fd_sc_hd__nor2_2 _21639_ (.A(_01836_),
    .B(_01837_),
    .Y(_01838_));
 sky130_fd_sc_hd__or2b_1 _21640_ (.A(_01693_),
    .B_N(_01698_),
    .X(_01839_));
 sky130_fd_sc_hd__or2b_1 _21641_ (.A(_01692_),
    .B_N(_01699_),
    .X(_01840_));
 sky130_fd_sc_hd__nand2_2 _21642_ (.A(_01839_),
    .B(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__and2b_1 _21643_ (.A_N(_01726_),
    .B(_01725_),
    .X(_01842_));
 sky130_fd_sc_hd__o21ba_1 _21644_ (.A1(_01694_),
    .A2(_01697_),
    .B1_N(_01695_),
    .X(_01843_));
 sky130_fd_sc_hd__buf_2 _21645_ (.A(_13836_),
    .X(_01844_));
 sky130_fd_sc_hd__a31o_1 _21646_ (.A1(_10894_),
    .A2(_01844_),
    .A3(_01716_),
    .B1(_01715_),
    .X(_01845_));
 sky130_fd_sc_hd__clkbuf_2 _21647_ (.A(_13605_),
    .X(_01846_));
 sky130_fd_sc_hd__a22oi_2 _21648_ (.A1(_13858_),
    .A2(_01846_),
    .B1(_13830_),
    .B2(_10784_),
    .Y(_01847_));
 sky130_fd_sc_hd__and4_1 _21649_ (.A(_13863_),
    .B(_14055_),
    .C(_13609_),
    .D(_14398_),
    .X(_01848_));
 sky130_fd_sc_hd__nor2_1 _21650_ (.A(_01847_),
    .B(_01848_),
    .Y(_01849_));
 sky130_fd_sc_hd__nand2_4 _21651_ (.A(\genblk1.pcpi_mul.rs2[6] ),
    .B(\genblk1.pcpi_mul.rs1[32] ),
    .Y(_01850_));
 sky130_fd_sc_hd__xnor2_1 _21652_ (.A(_01849_),
    .B(_01850_),
    .Y(_01851_));
 sky130_fd_sc_hd__xor2_1 _21653_ (.A(_01845_),
    .B(_01851_),
    .X(_01852_));
 sky130_fd_sc_hd__xnor2_1 _21654_ (.A(_01843_),
    .B(_01852_),
    .Y(_01853_));
 sky130_fd_sc_hd__o21ai_2 _21655_ (.A1(_01842_),
    .A2(_01728_),
    .B1(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__or3_1 _21656_ (.A(_01842_),
    .B(_01728_),
    .C(_01853_),
    .X(_01855_));
 sky130_fd_sc_hd__nand3_2 _21657_ (.A(_01841_),
    .B(_01854_),
    .C(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__a21o_1 _21658_ (.A1(_01854_),
    .A2(_01855_),
    .B1(_01841_),
    .X(_01857_));
 sky130_fd_sc_hd__nand2_1 _21659_ (.A(_01856_),
    .B(_01857_),
    .Y(_01858_));
 sky130_fd_sc_hd__nand2_2 _21660_ (.A(_01701_),
    .B(_01703_),
    .Y(_01859_));
 sky130_fd_sc_hd__xnor2_2 _21661_ (.A(_01858_),
    .B(_01859_),
    .Y(_01860_));
 sky130_fd_sc_hd__xnor2_1 _21662_ (.A(_01838_),
    .B(_01860_),
    .Y(_01861_));
 sky130_fd_sc_hd__xor2_2 _21663_ (.A(_01833_),
    .B(_01861_),
    .X(_01862_));
 sky130_fd_sc_hd__xor2_2 _21664_ (.A(_01832_),
    .B(_01862_),
    .X(_01863_));
 sky130_fd_sc_hd__nor2_1 _21665_ (.A(_01742_),
    .B(_01744_),
    .Y(_01864_));
 sky130_fd_sc_hd__a21o_1 _21666_ (.A1(_01752_),
    .A2(_01608_),
    .B1(_01768_),
    .X(_01865_));
 sky130_fd_sc_hd__buf_2 _21667_ (.A(_13838_),
    .X(_01866_));
 sky130_fd_sc_hd__a22oi_2 _21668_ (.A1(_13665_),
    .A2(_01866_),
    .B1(_13612_),
    .B2(_13670_),
    .Y(_01867_));
 sky130_fd_sc_hd__and4_1 _21669_ (.A(_13661_),
    .B(_13662_),
    .C(_13446_),
    .D(_01516_),
    .X(_01868_));
 sky130_fd_sc_hd__nor2_1 _21670_ (.A(_01867_),
    .B(_01868_),
    .Y(_01869_));
 sky130_fd_sc_hd__clkbuf_2 _21671_ (.A(_13813_),
    .X(_01870_));
 sky130_fd_sc_hd__nand2_1 _21672_ (.A(_11138_),
    .B(_01870_),
    .Y(_01871_));
 sky130_fd_sc_hd__xnor2_1 _21673_ (.A(_01869_),
    .B(_01871_),
    .Y(_01872_));
 sky130_fd_sc_hd__nand2_1 _21674_ (.A(_13897_),
    .B(_01538_),
    .Y(_01873_));
 sky130_fd_sc_hd__and4_1 _21675_ (.A(_11236_),
    .B(_13676_),
    .C(_12546_),
    .D(_13636_),
    .X(_01874_));
 sky130_fd_sc_hd__a22o_1 _21676_ (.A1(_14087_),
    .A2(_12546_),
    .B1(_13636_),
    .B2(_14086_),
    .X(_01875_));
 sky130_fd_sc_hd__and2b_1 _21677_ (.A_N(_01874_),
    .B(_01875_),
    .X(_01876_));
 sky130_fd_sc_hd__xnor2_1 _21678_ (.A(_01873_),
    .B(_01876_),
    .Y(_01877_));
 sky130_fd_sc_hd__o21ba_1 _21679_ (.A1(_01721_),
    .A2(_01723_),
    .B1_N(_01722_),
    .X(_01878_));
 sky130_fd_sc_hd__xnor2_1 _21680_ (.A(_01877_),
    .B(_01878_),
    .Y(_01879_));
 sky130_fd_sc_hd__and2_1 _21681_ (.A(_01872_),
    .B(_01879_),
    .X(_01880_));
 sky130_fd_sc_hd__nor2_1 _21682_ (.A(_01872_),
    .B(_01879_),
    .Y(_01881_));
 sky130_fd_sc_hd__or2_2 _21683_ (.A(_01880_),
    .B(_01881_),
    .X(_01882_));
 sky130_fd_sc_hd__or2b_1 _21684_ (.A(_01734_),
    .B_N(_01739_),
    .X(_01883_));
 sky130_fd_sc_hd__nand2_1 _21685_ (.A(_01733_),
    .B(_01740_),
    .Y(_01884_));
 sky130_fd_sc_hd__clkbuf_2 _21686_ (.A(_13891_),
    .X(_01885_));
 sky130_fd_sc_hd__a31o_1 _21687_ (.A1(_14099_),
    .A2(_01885_),
    .A3(_01737_),
    .B1(_01736_),
    .X(_01886_));
 sky130_fd_sc_hd__o21ba_1 _21688_ (.A1(_01753_),
    .A2(_01758_),
    .B1_N(_01756_),
    .X(_01887_));
 sky130_fd_sc_hd__a22oi_1 _21689_ (.A1(_11782_),
    .A2(_13484_),
    .B1(_12694_),
    .B2(_11664_),
    .Y(_01888_));
 sky130_fd_sc_hd__and4_1 _21690_ (.A(_11656_),
    .B(_11659_),
    .C(_12274_),
    .D(_14268_),
    .X(_01889_));
 sky130_fd_sc_hd__nor2_1 _21691_ (.A(_01888_),
    .B(_01889_),
    .Y(_01890_));
 sky130_fd_sc_hd__nand2_1 _21692_ (.A(_11445_),
    .B(_13888_),
    .Y(_01891_));
 sky130_fd_sc_hd__xnor2_2 _21693_ (.A(_01890_),
    .B(_01891_),
    .Y(_01892_));
 sky130_fd_sc_hd__xnor2_1 _21694_ (.A(_01887_),
    .B(_01892_),
    .Y(_01893_));
 sky130_fd_sc_hd__xnor2_1 _21695_ (.A(_01886_),
    .B(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__a21oi_1 _21696_ (.A1(_01883_),
    .A2(_01884_),
    .B1(_01894_),
    .Y(_01895_));
 sky130_fd_sc_hd__and3_1 _21697_ (.A(_01883_),
    .B(_01884_),
    .C(_01894_),
    .X(_01896_));
 sky130_fd_sc_hd__nor3_1 _21698_ (.A(_01882_),
    .B(_01895_),
    .C(_01896_),
    .Y(_01897_));
 sky130_fd_sc_hd__o21a_1 _21699_ (.A1(_01895_),
    .A2(_01896_),
    .B1(_01882_),
    .X(_01898_));
 sky130_fd_sc_hd__a211oi_1 _21700_ (.A1(_01865_),
    .A2(_01771_),
    .B1(_01897_),
    .C1(_01898_),
    .Y(_01899_));
 sky130_fd_sc_hd__o211ai_1 _21701_ (.A1(_01897_),
    .A2(_01898_),
    .B1(_01865_),
    .C1(_01771_),
    .Y(_01900_));
 sky130_fd_sc_hd__and2b_1 _21702_ (.A_N(_01899_),
    .B(_01900_),
    .X(_01901_));
 sky130_fd_sc_hd__xnor2_2 _21703_ (.A(_01864_),
    .B(_01901_),
    .Y(_01902_));
 sky130_fd_sc_hd__or2b_1 _21704_ (.A(_01766_),
    .B_N(_01765_),
    .X(_01903_));
 sky130_fd_sc_hd__nand2_1 _21705_ (.A(_01760_),
    .B(_01767_),
    .Y(_01904_));
 sky130_fd_sc_hd__or3_1 _21706_ (.A(_01774_),
    .B(_01777_),
    .C(_01778_),
    .X(_01905_));
 sky130_fd_sc_hd__nand2_1 _21707_ (.A(_12591_),
    .B(_13663_),
    .Y(_01906_));
 sky130_fd_sc_hd__and4_1 _21708_ (.A(_13679_),
    .B(_13713_),
    .C(_11959_),
    .D(_13715_),
    .X(_01907_));
 sky130_fd_sc_hd__a22oi_1 _21709_ (.A1(_11896_),
    .A2(_13901_),
    .B1(_13716_),
    .B2(_11950_),
    .Y(_01908_));
 sky130_fd_sc_hd__nor2_1 _21710_ (.A(_01907_),
    .B(_01908_),
    .Y(_01909_));
 sky130_fd_sc_hd__xnor2_2 _21711_ (.A(_01906_),
    .B(_01909_),
    .Y(_01910_));
 sky130_fd_sc_hd__nand2_1 _21712_ (.A(_12075_),
    .B(_12227_),
    .Y(_01911_));
 sky130_fd_sc_hd__clkbuf_2 _21713_ (.A(_12322_),
    .X(_01912_));
 sky130_fd_sc_hd__and4_1 _21714_ (.A(_11490_),
    .B(_13689_),
    .C(_01912_),
    .D(_13944_),
    .X(_01913_));
 sky130_fd_sc_hd__a22oi_2 _21715_ (.A1(_11599_),
    .A2(_13942_),
    .B1(_13721_),
    .B2(_11825_),
    .Y(_01914_));
 sky130_fd_sc_hd__nor2_1 _21716_ (.A(_01913_),
    .B(_01914_),
    .Y(_01915_));
 sky130_fd_sc_hd__xnor2_1 _21717_ (.A(_01911_),
    .B(_01915_),
    .Y(_01916_));
 sky130_fd_sc_hd__o21ba_1 _21718_ (.A1(_01761_),
    .A2(_01763_),
    .B1_N(_01762_),
    .X(_01917_));
 sky130_fd_sc_hd__xnor2_1 _21719_ (.A(_01916_),
    .B(_01917_),
    .Y(_01918_));
 sky130_fd_sc_hd__xnor2_1 _21720_ (.A(_01910_),
    .B(_01918_),
    .Y(_01919_));
 sky130_fd_sc_hd__a21oi_1 _21721_ (.A1(_01905_),
    .A2(_01781_),
    .B1(_01919_),
    .Y(_01920_));
 sky130_fd_sc_hd__and3_1 _21722_ (.A(_01905_),
    .B(_01781_),
    .C(_01919_),
    .X(_01921_));
 sky130_fd_sc_hd__a211o_1 _21723_ (.A1(_01903_),
    .A2(_01904_),
    .B1(_01920_),
    .C1(_01921_),
    .X(_01922_));
 sky130_fd_sc_hd__o211ai_1 _21724_ (.A1(_01920_),
    .A2(_01921_),
    .B1(_01903_),
    .C1(_01904_),
    .Y(_01923_));
 sky130_fd_sc_hd__and2_1 _21725_ (.A(_01922_),
    .B(_01923_),
    .X(_01924_));
 sky130_fd_sc_hd__o21ba_1 _21726_ (.A1(_01784_),
    .A2(_01786_),
    .B1_N(_01785_),
    .X(_01925_));
 sky130_fd_sc_hd__and4_1 _21727_ (.A(_11601_),
    .B(_11372_),
    .C(_13555_),
    .D(_13556_),
    .X(_01926_));
 sky130_fd_sc_hd__a22oi_2 _21728_ (.A1(_12343_),
    .A2(_13743_),
    .B1(_13744_),
    .B2(_11473_),
    .Y(_01927_));
 sky130_fd_sc_hd__and4bb_1 _21729_ (.A_N(_01926_),
    .B_N(_01927_),
    .C(_11477_),
    .D(_12585_),
    .X(_01928_));
 sky130_fd_sc_hd__o2bb2a_1 _21730_ (.A1_N(_11477_),
    .A2_N(_14147_),
    .B1(_01926_),
    .B2(_01927_),
    .X(_01929_));
 sky130_fd_sc_hd__nor2_1 _21731_ (.A(_01928_),
    .B(_01929_),
    .Y(_01930_));
 sky130_fd_sc_hd__xnor2_1 _21732_ (.A(_01925_),
    .B(_01930_),
    .Y(_01931_));
 sky130_fd_sc_hd__o21ai_2 _21733_ (.A1(_01775_),
    .A2(_01777_),
    .B1(_01931_),
    .Y(_01932_));
 sky130_fd_sc_hd__or3_1 _21734_ (.A(_01775_),
    .B(_01777_),
    .C(_01931_),
    .X(_01933_));
 sky130_fd_sc_hd__and2_1 _21735_ (.A(_01932_),
    .B(_01933_),
    .X(_01934_));
 sky130_fd_sc_hd__nand2_1 _21736_ (.A(_11161_),
    .B(_13226_),
    .Y(_01935_));
 sky130_fd_sc_hd__and4_1 _21737_ (.A(_11037_),
    .B(_11043_),
    .C(_13228_),
    .D(_14508_),
    .X(_01936_));
 sky130_fd_sc_hd__a22oi_1 _21738_ (.A1(_11270_),
    .A2(_13970_),
    .B1(_14510_),
    .B2(_11386_),
    .Y(_01937_));
 sky130_fd_sc_hd__nor2_1 _21739_ (.A(_01936_),
    .B(_01937_),
    .Y(_01938_));
 sky130_fd_sc_hd__xnor2_2 _21740_ (.A(_01935_),
    .B(_01938_),
    .Y(_01939_));
 sky130_fd_sc_hd__nand2_1 _21741_ (.A(_11402_),
    .B(_14160_),
    .Y(_01940_));
 sky130_fd_sc_hd__and2b_1 _21742_ (.A_N(_10757_),
    .B(_01618_),
    .X(_01941_));
 sky130_fd_sc_hd__nand2_1 _21743_ (.A(_11059_),
    .B(_13753_),
    .Y(_01942_));
 sky130_fd_sc_hd__xnor2_1 _21744_ (.A(_01941_),
    .B(_01942_),
    .Y(_01943_));
 sky130_fd_sc_hd__xnor2_1 _21745_ (.A(_01940_),
    .B(_01943_),
    .Y(_01944_));
 sky130_fd_sc_hd__and3_1 _21746_ (.A(_11404_),
    .B(_13757_),
    .C(_01790_),
    .X(_01945_));
 sky130_fd_sc_hd__a31o_1 _21747_ (.A1(_11297_),
    .A2(_14166_),
    .A3(_01792_),
    .B1(_01945_),
    .X(_01946_));
 sky130_fd_sc_hd__xor2_1 _21748_ (.A(_01944_),
    .B(_01946_),
    .X(_01947_));
 sky130_fd_sc_hd__xnor2_1 _21749_ (.A(_01939_),
    .B(_01947_),
    .Y(_01948_));
 sky130_fd_sc_hd__nand2_1 _21750_ (.A(_01793_),
    .B(_01795_),
    .Y(_01949_));
 sky130_fd_sc_hd__a21boi_1 _21751_ (.A1(_01788_),
    .A2(_01796_),
    .B1_N(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__xnor2_1 _21752_ (.A(_01948_),
    .B(_01950_),
    .Y(_01951_));
 sky130_fd_sc_hd__xnor2_2 _21753_ (.A(_01934_),
    .B(_01951_),
    .Y(_01952_));
 sky130_fd_sc_hd__nand2_1 _21754_ (.A(_01797_),
    .B(_01799_),
    .Y(_01953_));
 sky130_fd_sc_hd__nor2_1 _21755_ (.A(_01797_),
    .B(_01799_),
    .Y(_01954_));
 sky130_fd_sc_hd__a21oi_2 _21756_ (.A1(_01783_),
    .A2(_01953_),
    .B1(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__xnor2_2 _21757_ (.A(_01952_),
    .B(_01955_),
    .Y(_01956_));
 sky130_fd_sc_hd__xnor2_2 _21758_ (.A(_01924_),
    .B(_01956_),
    .Y(_01957_));
 sky130_fd_sc_hd__and2b_1 _21759_ (.A_N(_01804_),
    .B(_01801_),
    .X(_01958_));
 sky130_fd_sc_hd__a21oi_2 _21760_ (.A1(_01773_),
    .A2(_01805_),
    .B1(_01958_),
    .Y(_01959_));
 sky130_fd_sc_hd__xor2_2 _21761_ (.A(_01957_),
    .B(_01959_),
    .X(_01960_));
 sky130_fd_sc_hd__xor2_2 _21762_ (.A(_01902_),
    .B(_01960_),
    .X(_01961_));
 sky130_fd_sc_hd__nor2_1 _21763_ (.A(_01806_),
    .B(_01808_),
    .Y(_01962_));
 sky130_fd_sc_hd__a21oi_2 _21764_ (.A1(_01749_),
    .A2(_01809_),
    .B1(_01962_),
    .Y(_01963_));
 sky130_fd_sc_hd__xnor2_2 _21765_ (.A(_01961_),
    .B(_01963_),
    .Y(_01964_));
 sky130_fd_sc_hd__xnor2_2 _21766_ (.A(_01863_),
    .B(_01964_),
    .Y(_01965_));
 sky130_fd_sc_hd__and2b_1 _21767_ (.A_N(_01812_),
    .B(_01810_),
    .X(_01966_));
 sky130_fd_sc_hd__a21oi_2 _21768_ (.A1(_01710_),
    .A2(_01813_),
    .B1(_01966_),
    .Y(_01967_));
 sky130_fd_sc_hd__xnor2_4 _21769_ (.A(_01965_),
    .B(_01967_),
    .Y(_01968_));
 sky130_fd_sc_hd__xnor2_4 _21770_ (.A(_01831_),
    .B(_01968_),
    .Y(_01969_));
 sky130_fd_sc_hd__or2b_1 _21771_ (.A(_01816_),
    .B_N(_01814_),
    .X(_01970_));
 sky130_fd_sc_hd__a21boi_4 _21772_ (.A1(_01674_),
    .A2(_01817_),
    .B1_N(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hd__xor2_4 _21773_ (.A(_01969_),
    .B(_01971_),
    .X(_01972_));
 sky130_fd_sc_hd__xnor2_4 _21774_ (.A(_01672_),
    .B(_01972_),
    .Y(_01973_));
 sky130_fd_sc_hd__nor2_1 _21775_ (.A(_01818_),
    .B(_01820_),
    .Y(_01974_));
 sky130_fd_sc_hd__a21oi_2 _21776_ (.A1(_14555_),
    .A2(_01821_),
    .B1(_01974_),
    .Y(_01975_));
 sky130_fd_sc_hd__xor2_4 _21777_ (.A(_01973_),
    .B(_01975_),
    .X(_01976_));
 sky130_fd_sc_hd__nand2_1 _21778_ (.A(_01657_),
    .B(_01823_),
    .Y(_01977_));
 sky130_fd_sc_hd__and3b_1 _21779_ (.A_N(_01659_),
    .B(_01666_),
    .C(_01825_),
    .X(_01978_));
 sky130_fd_sc_hd__a21oi_2 _21780_ (.A1(_01824_),
    .A2(_01977_),
    .B1(_01978_),
    .Y(_01979_));
 sky130_fd_sc_hd__xnor2_4 _21781_ (.A(_01976_),
    .B(_01979_),
    .Y(_00084_));
 sky130_fd_sc_hd__nor2_1 _21782_ (.A(_01969_),
    .B(_01971_),
    .Y(_01980_));
 sky130_fd_sc_hd__a21oi_4 _21783_ (.A1(_01672_),
    .A2(_01972_),
    .B1(_01980_),
    .Y(_01981_));
 sky130_fd_sc_hd__nor2_2 _21784_ (.A(_01829_),
    .B(_01830_),
    .Y(_01982_));
 sky130_fd_sc_hd__nand2_1 _21785_ (.A(_01838_),
    .B(_01860_),
    .Y(_01983_));
 sky130_fd_sc_hd__or2_1 _21786_ (.A(_01838_),
    .B(_01860_),
    .X(_01984_));
 sky130_fd_sc_hd__nor2_1 _21787_ (.A(_01832_),
    .B(_01862_),
    .Y(_01985_));
 sky130_fd_sc_hd__a31o_1 _21788_ (.A1(_01833_),
    .A2(_01983_),
    .A3(_01984_),
    .B1(_01985_),
    .X(_01986_));
 sky130_fd_sc_hd__and3_2 _21789_ (.A(_10586_),
    .B(_14396_),
    .C(_01678_),
    .X(_01987_));
 sky130_fd_sc_hd__nor2_1 _21790_ (.A(_01987_),
    .B(_01836_),
    .Y(_01988_));
 sky130_fd_sc_hd__xnor2_2 _21791_ (.A(_01986_),
    .B(_01988_),
    .Y(_01989_));
 sky130_fd_sc_hd__a32oi_4 _21792_ (.A1(_01856_),
    .A2(_01857_),
    .A3(_01859_),
    .B1(_01860_),
    .B2(_01838_),
    .Y(_01990_));
 sky130_fd_sc_hd__or3b_1 _21793_ (.A(_01864_),
    .B(_01899_),
    .C_N(_01900_),
    .X(_01991_));
 sky130_fd_sc_hd__and2b_1 _21794_ (.A_N(_01899_),
    .B(_01991_),
    .X(_01992_));
 sky130_fd_sc_hd__o21ba_1 _21795_ (.A1(_14396_),
    .A2(_01834_),
    .B1_N(_01987_),
    .X(_01993_));
 sky130_fd_sc_hd__xnor2_1 _21796_ (.A(_14566_),
    .B(_01993_),
    .Y(_01994_));
 sky130_fd_sc_hd__clkbuf_4 _21797_ (.A(_01994_),
    .X(_01995_));
 sky130_fd_sc_hd__or2b_1 _21798_ (.A(_01843_),
    .B_N(_01852_),
    .X(_01996_));
 sky130_fd_sc_hd__a21bo_1 _21799_ (.A1(_01845_),
    .A2(_01851_),
    .B1_N(_01996_),
    .X(_01997_));
 sky130_fd_sc_hd__and2b_1 _21800_ (.A_N(_01878_),
    .B(_01877_),
    .X(_01998_));
 sky130_fd_sc_hd__o21ba_1 _21801_ (.A1(_01847_),
    .A2(_01850_),
    .B1_N(_01848_),
    .X(_01999_));
 sky130_fd_sc_hd__o21ba_1 _21802_ (.A1(_01867_),
    .A2(_01871_),
    .B1_N(_01868_),
    .X(_02000_));
 sky130_fd_sc_hd__and3_4 _21803_ (.A(_10781_),
    .B(\genblk1.pcpi_mul.rs2[8] ),
    .C(\genblk1.pcpi_mul.rs1[32] ),
    .X(_02001_));
 sky130_fd_sc_hd__a22o_1 _21804_ (.A1(_11201_),
    .A2(\genblk1.pcpi_mul.rs1[31] ),
    .B1(_14024_),
    .B2(_10783_),
    .X(_02002_));
 sky130_fd_sc_hd__a21bo_1 _21805_ (.A1(_14210_),
    .A2(_02001_),
    .B1_N(_02002_),
    .X(_02003_));
 sky130_fd_sc_hd__xor2_1 _21806_ (.A(_01850_),
    .B(_02003_),
    .X(_02004_));
 sky130_fd_sc_hd__xnor2_1 _21807_ (.A(_02000_),
    .B(_02004_),
    .Y(_02005_));
 sky130_fd_sc_hd__xnor2_1 _21808_ (.A(_01999_),
    .B(_02005_),
    .Y(_02006_));
 sky130_fd_sc_hd__o21ai_1 _21809_ (.A1(_01998_),
    .A2(_01880_),
    .B1(_02006_),
    .Y(_02007_));
 sky130_fd_sc_hd__or3_1 _21810_ (.A(_01998_),
    .B(_01880_),
    .C(_02006_),
    .X(_02008_));
 sky130_fd_sc_hd__and3_1 _21811_ (.A(_01997_),
    .B(_02007_),
    .C(_02008_),
    .X(_02009_));
 sky130_fd_sc_hd__a21oi_1 _21812_ (.A1(_02007_),
    .A2(_02008_),
    .B1(_01997_),
    .Y(_02010_));
 sky130_fd_sc_hd__nor2_1 _21813_ (.A(_02009_),
    .B(_02010_),
    .Y(_02011_));
 sky130_fd_sc_hd__nand2_1 _21814_ (.A(_01854_),
    .B(_01856_),
    .Y(_02012_));
 sky130_fd_sc_hd__xnor2_1 _21815_ (.A(_02011_),
    .B(_02012_),
    .Y(_02013_));
 sky130_fd_sc_hd__xor2_1 _21816_ (.A(_01995_),
    .B(_02013_),
    .X(_02014_));
 sky130_fd_sc_hd__xnor2_1 _21817_ (.A(_01992_),
    .B(_02014_),
    .Y(_02015_));
 sky130_fd_sc_hd__xnor2_2 _21818_ (.A(_01990_),
    .B(_02015_),
    .Y(_02016_));
 sky130_fd_sc_hd__nor2_1 _21819_ (.A(_01895_),
    .B(_01897_),
    .Y(_02017_));
 sky130_fd_sc_hd__a21o_1 _21820_ (.A1(_01905_),
    .A2(_01781_),
    .B1(_01919_),
    .X(_02018_));
 sky130_fd_sc_hd__a22o_1 _21821_ (.A1(_11145_),
    .A2(_13281_),
    .B1(_13608_),
    .B2(_10957_),
    .X(_02019_));
 sky130_fd_sc_hd__nand4_1 _21822_ (.A(_13669_),
    .B(_11108_),
    .C(_14418_),
    .D(_13608_),
    .Y(_02020_));
 sky130_fd_sc_hd__and2_1 _21823_ (.A(_11900_),
    .B(_13605_),
    .X(_02021_));
 sky130_fd_sc_hd__a21oi_1 _21824_ (.A1(_02019_),
    .A2(_02020_),
    .B1(_02021_),
    .Y(_02022_));
 sky130_fd_sc_hd__and3_2 _21825_ (.A(_02019_),
    .B(_02020_),
    .C(_02021_),
    .X(_02023_));
 sky130_fd_sc_hd__nor2_1 _21826_ (.A(_02022_),
    .B(_02023_),
    .Y(_02024_));
 sky130_fd_sc_hd__nand2_1 _21827_ (.A(_11135_),
    .B(_14417_),
    .Y(_02025_));
 sky130_fd_sc_hd__nand4_1 _21828_ (.A(_13680_),
    .B(_13678_),
    .C(_13125_),
    .D(_13285_),
    .Y(_02026_));
 sky130_fd_sc_hd__a22o_1 _21829_ (.A1(_13678_),
    .A2(_13632_),
    .B1(_13285_),
    .B2(_14086_),
    .X(_02027_));
 sky130_fd_sc_hd__nand3b_1 _21830_ (.A_N(_02025_),
    .B(_02026_),
    .C(_02027_),
    .Y(_02028_));
 sky130_fd_sc_hd__a21bo_1 _21831_ (.A1(_02026_),
    .A2(_02027_),
    .B1_N(_02025_),
    .X(_02029_));
 sky130_fd_sc_hd__nand2_1 _21832_ (.A(_02028_),
    .B(_02029_),
    .Y(_02030_));
 sky130_fd_sc_hd__a31o_1 _21833_ (.A1(_11233_),
    .A2(_14438_),
    .A3(_01875_),
    .B1(_01874_),
    .X(_02031_));
 sky130_fd_sc_hd__xnor2_2 _21834_ (.A(_02030_),
    .B(_02031_),
    .Y(_02032_));
 sky130_fd_sc_hd__xnor2_2 _21835_ (.A(_02024_),
    .B(_02032_),
    .Y(_02033_));
 sky130_fd_sc_hd__or2b_1 _21836_ (.A(_01887_),
    .B_N(_01892_),
    .X(_02034_));
 sky130_fd_sc_hd__nand2_1 _21837_ (.A(_01886_),
    .B(_01893_),
    .Y(_02035_));
 sky130_fd_sc_hd__buf_2 _21838_ (.A(_13888_),
    .X(_02036_));
 sky130_fd_sc_hd__a31o_1 _21839_ (.A1(_11446_),
    .A2(_02036_),
    .A3(_01890_),
    .B1(_01889_),
    .X(_02037_));
 sky130_fd_sc_hd__o21ba_1 _21840_ (.A1(_01906_),
    .A2(_01908_),
    .B1_N(_01907_),
    .X(_02038_));
 sky130_fd_sc_hd__a22oi_1 _21841_ (.A1(_11665_),
    .A2(_12282_),
    .B1(_12830_),
    .B2(_14103_),
    .Y(_02039_));
 sky130_fd_sc_hd__and4_1 _21842_ (.A(_11923_),
    .B(_11781_),
    .C(_12983_),
    .D(_12538_),
    .X(_02040_));
 sky130_fd_sc_hd__nor2_1 _21843_ (.A(_02039_),
    .B(_02040_),
    .Y(_02041_));
 sky130_fd_sc_hd__nand2_1 _21844_ (.A(_11444_),
    .B(_12977_),
    .Y(_02042_));
 sky130_fd_sc_hd__xnor2_2 _21845_ (.A(_02041_),
    .B(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__xnor2_1 _21846_ (.A(_02038_),
    .B(_02043_),
    .Y(_02044_));
 sky130_fd_sc_hd__xnor2_1 _21847_ (.A(_02037_),
    .B(_02044_),
    .Y(_02045_));
 sky130_fd_sc_hd__a21oi_1 _21848_ (.A1(_02034_),
    .A2(_02035_),
    .B1(_02045_),
    .Y(_02046_));
 sky130_fd_sc_hd__and3_1 _21849_ (.A(_02034_),
    .B(_02035_),
    .C(_02045_),
    .X(_02047_));
 sky130_fd_sc_hd__nor3_1 _21850_ (.A(_02033_),
    .B(_02046_),
    .C(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__o21a_1 _21851_ (.A1(_02046_),
    .A2(_02047_),
    .B1(_02033_),
    .X(_02049_));
 sky130_fd_sc_hd__a211oi_1 _21852_ (.A1(_02018_),
    .A2(_01922_),
    .B1(net355),
    .C1(_02049_),
    .Y(_02050_));
 sky130_fd_sc_hd__o211ai_1 _21853_ (.A1(net355),
    .A2(_02049_),
    .B1(_02018_),
    .C1(_01922_),
    .Y(_02051_));
 sky130_fd_sc_hd__and2b_1 _21854_ (.A_N(_02050_),
    .B(_02051_),
    .X(_02052_));
 sky130_fd_sc_hd__xnor2_2 _21855_ (.A(_02017_),
    .B(_02052_),
    .Y(_02053_));
 sky130_fd_sc_hd__or2b_1 _21856_ (.A(_01917_),
    .B_N(_01916_),
    .X(_02054_));
 sky130_fd_sc_hd__nand2_1 _21857_ (.A(_01910_),
    .B(_01918_),
    .Y(_02055_));
 sky130_fd_sc_hd__or3_1 _21858_ (.A(_01925_),
    .B(_01928_),
    .C(_01929_),
    .X(_02056_));
 sky130_fd_sc_hd__nand2_1 _21859_ (.A(_11770_),
    .B(_12274_),
    .Y(_02057_));
 sky130_fd_sc_hd__and4_1 _21860_ (.A(_11890_),
    .B(_13305_),
    .C(_12021_),
    .D(_12079_),
    .X(_02058_));
 sky130_fd_sc_hd__a22oi_1 _21861_ (.A1(_11959_),
    .A2(_13715_),
    .B1(_12145_),
    .B2(_13713_),
    .Y(_02059_));
 sky130_fd_sc_hd__nor2_1 _21862_ (.A(_02058_),
    .B(_02059_),
    .Y(_02060_));
 sky130_fd_sc_hd__xnor2_2 _21863_ (.A(_02057_),
    .B(_02060_),
    .Y(_02061_));
 sky130_fd_sc_hd__nand2_1 _21864_ (.A(_11950_),
    .B(_14482_),
    .Y(_02062_));
 sky130_fd_sc_hd__and4_1 _21865_ (.A(_13689_),
    .B(_12074_),
    .C(_01912_),
    .D(_13944_),
    .X(_02063_));
 sky130_fd_sc_hd__a22oi_2 _21866_ (.A1(_13918_),
    .A2(_12329_),
    .B1(_13721_),
    .B2(_11599_),
    .Y(_02064_));
 sky130_fd_sc_hd__nor2_1 _21867_ (.A(_02063_),
    .B(_02064_),
    .Y(_02065_));
 sky130_fd_sc_hd__xnor2_1 _21868_ (.A(_02062_),
    .B(_02065_),
    .Y(_02066_));
 sky130_fd_sc_hd__o21ba_1 _21869_ (.A1(_01911_),
    .A2(_01914_),
    .B1_N(_01913_),
    .X(_02067_));
 sky130_fd_sc_hd__xnor2_1 _21870_ (.A(_02066_),
    .B(_02067_),
    .Y(_02068_));
 sky130_fd_sc_hd__xnor2_1 _21871_ (.A(_02061_),
    .B(_02068_),
    .Y(_02069_));
 sky130_fd_sc_hd__a21oi_2 _21872_ (.A1(_02056_),
    .A2(_01932_),
    .B1(_02069_),
    .Y(_02070_));
 sky130_fd_sc_hd__and3_1 _21873_ (.A(_02056_),
    .B(_01932_),
    .C(_02069_),
    .X(_02071_));
 sky130_fd_sc_hd__a211oi_2 _21874_ (.A1(_02054_),
    .A2(_02055_),
    .B1(_02070_),
    .C1(_02071_),
    .Y(_02072_));
 sky130_fd_sc_hd__o211a_1 _21875_ (.A1(_02070_),
    .A2(_02071_),
    .B1(_02054_),
    .C1(_02055_),
    .X(_02073_));
 sky130_fd_sc_hd__nor2_2 _21876_ (.A(_02072_),
    .B(_02073_),
    .Y(_02074_));
 sky130_fd_sc_hd__o21ba_1 _21877_ (.A1(_01935_),
    .A2(_01937_),
    .B1_N(_01936_),
    .X(_02075_));
 sky130_fd_sc_hd__a22oi_1 _21878_ (.A1(_11482_),
    .A2(_13743_),
    .B1(_13744_),
    .B2(_11479_),
    .Y(_02076_));
 sky130_fd_sc_hd__and4_1 _21879_ (.A(_11277_),
    .B(_11380_),
    .C(_12776_),
    .D(_13556_),
    .X(_02077_));
 sky130_fd_sc_hd__o2bb2a_1 _21880_ (.A1_N(_11491_),
    .A2_N(_14147_),
    .B1(_02076_),
    .B2(_02077_),
    .X(_02078_));
 sky130_fd_sc_hd__and4bb_1 _21881_ (.A_N(_02076_),
    .B_N(_02077_),
    .C(_11491_),
    .D(_14147_),
    .X(_02079_));
 sky130_fd_sc_hd__nor2_1 _21882_ (.A(_02078_),
    .B(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__xnor2_1 _21883_ (.A(_02075_),
    .B(_02080_),
    .Y(_02081_));
 sky130_fd_sc_hd__o21ai_2 _21884_ (.A1(_01926_),
    .A2(_01928_),
    .B1(_02081_),
    .Y(_02082_));
 sky130_fd_sc_hd__or3_1 _21885_ (.A(_01926_),
    .B(_01928_),
    .C(_02081_),
    .X(_02083_));
 sky130_fd_sc_hd__and2_2 _21886_ (.A(_02082_),
    .B(_02083_),
    .X(_02084_));
 sky130_fd_sc_hd__nand2_1 _21887_ (.A(_11262_),
    .B(_13055_),
    .Y(_02085_));
 sky130_fd_sc_hd__and4_1 _21888_ (.A(_11156_),
    .B(_11264_),
    .C(_13764_),
    .D(_13765_),
    .X(_02086_));
 sky130_fd_sc_hd__a22oi_2 _21889_ (.A1(_11068_),
    .A2(_13970_),
    .B1(_13972_),
    .B2(_11270_),
    .Y(_02087_));
 sky130_fd_sc_hd__nor2_1 _21890_ (.A(_02086_),
    .B(_02087_),
    .Y(_02088_));
 sky130_fd_sc_hd__xnor2_2 _21891_ (.A(_02085_),
    .B(_02088_),
    .Y(_02089_));
 sky130_fd_sc_hd__nand2_1 _21892_ (.A(_11167_),
    .B(_14160_),
    .Y(_02090_));
 sky130_fd_sc_hd__and2b_1 _21893_ (.A_N(_10852_),
    .B(_13802_),
    .X(_02091_));
 sky130_fd_sc_hd__nand2_1 _21894_ (.A(_11175_),
    .B(_13756_),
    .Y(_02092_));
 sky130_fd_sc_hd__xnor2_2 _21895_ (.A(_02091_),
    .B(_02092_),
    .Y(_02093_));
 sky130_fd_sc_hd__xnor2_2 _21896_ (.A(_02090_),
    .B(_02093_),
    .Y(_02094_));
 sky130_fd_sc_hd__and3_1 _21897_ (.A(_13959_),
    .B(_13757_),
    .C(_01941_),
    .X(_02095_));
 sky130_fd_sc_hd__a31o_1 _21898_ (.A1(_11050_),
    .A2(_14166_),
    .A3(_01943_),
    .B1(_02095_),
    .X(_02096_));
 sky130_fd_sc_hd__xor2_2 _21899_ (.A(_02094_),
    .B(_02096_),
    .X(_02097_));
 sky130_fd_sc_hd__xnor2_2 _21900_ (.A(_02089_),
    .B(_02097_),
    .Y(_02098_));
 sky130_fd_sc_hd__nand2_1 _21901_ (.A(_01944_),
    .B(_01946_),
    .Y(_02099_));
 sky130_fd_sc_hd__a21boi_2 _21902_ (.A1(_01939_),
    .A2(_01947_),
    .B1_N(_02099_),
    .Y(_02100_));
 sky130_fd_sc_hd__xnor2_2 _21903_ (.A(_02098_),
    .B(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__xnor2_4 _21904_ (.A(_02084_),
    .B(_02101_),
    .Y(_02102_));
 sky130_fd_sc_hd__nand2_1 _21905_ (.A(_01948_),
    .B(_01950_),
    .Y(_02103_));
 sky130_fd_sc_hd__nor2_1 _21906_ (.A(_01948_),
    .B(_01950_),
    .Y(_02104_));
 sky130_fd_sc_hd__a21oi_2 _21907_ (.A1(_01934_),
    .A2(_02103_),
    .B1(_02104_),
    .Y(_02105_));
 sky130_fd_sc_hd__xnor2_4 _21908_ (.A(_02102_),
    .B(_02105_),
    .Y(_02106_));
 sky130_fd_sc_hd__xnor2_2 _21909_ (.A(_02074_),
    .B(_02106_),
    .Y(_02107_));
 sky130_fd_sc_hd__and2b_1 _21910_ (.A_N(_01955_),
    .B(_01952_),
    .X(_02108_));
 sky130_fd_sc_hd__a21oi_2 _21911_ (.A1(_01924_),
    .A2(_01956_),
    .B1(_02108_),
    .Y(_02109_));
 sky130_fd_sc_hd__xor2_2 _21912_ (.A(_02107_),
    .B(_02109_),
    .X(_02110_));
 sky130_fd_sc_hd__xor2_2 _21913_ (.A(_02053_),
    .B(_02110_),
    .X(_02111_));
 sky130_fd_sc_hd__nor2_1 _21914_ (.A(_01957_),
    .B(_01959_),
    .Y(_02112_));
 sky130_fd_sc_hd__a21oi_2 _21915_ (.A1(_01902_),
    .A2(_01960_),
    .B1(_02112_),
    .Y(_02113_));
 sky130_fd_sc_hd__xnor2_2 _21916_ (.A(_02111_),
    .B(_02113_),
    .Y(_02114_));
 sky130_fd_sc_hd__xnor2_2 _21917_ (.A(_02016_),
    .B(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__or2b_1 _21918_ (.A(_01963_),
    .B_N(_01961_),
    .X(_02116_));
 sky130_fd_sc_hd__a21boi_2 _21919_ (.A1(_01863_),
    .A2(_01964_),
    .B1_N(_02116_),
    .Y(_02117_));
 sky130_fd_sc_hd__xor2_2 _21920_ (.A(_02115_),
    .B(_02117_),
    .X(_02118_));
 sky130_fd_sc_hd__xor2_2 _21921_ (.A(_01989_),
    .B(_02118_),
    .X(_02119_));
 sky130_fd_sc_hd__or2_1 _21922_ (.A(_01965_),
    .B(_01967_),
    .X(_02120_));
 sky130_fd_sc_hd__o21a_1 _21923_ (.A1(_01831_),
    .A2(_01968_),
    .B1(_02120_),
    .X(_02121_));
 sky130_fd_sc_hd__xnor2_2 _21924_ (.A(_02119_),
    .B(_02121_),
    .Y(_02122_));
 sky130_fd_sc_hd__xnor2_4 _21925_ (.A(_01982_),
    .B(_02122_),
    .Y(_02123_));
 sky130_fd_sc_hd__xor2_4 _21926_ (.A(_01981_),
    .B(_02123_),
    .X(_02124_));
 sky130_fd_sc_hd__or2_1 _21927_ (.A(_01973_),
    .B(_01975_),
    .X(_02125_));
 sky130_fd_sc_hd__or2b_1 _21928_ (.A(_01979_),
    .B_N(_01976_),
    .X(_02126_));
 sky130_fd_sc_hd__nand2_2 _21929_ (.A(_02125_),
    .B(_02126_),
    .Y(_02127_));
 sky130_fd_sc_hd__xor2_4 _21930_ (.A(_02124_),
    .B(_02127_),
    .X(_00085_));
 sky130_fd_sc_hd__o21a_1 _21931_ (.A1(_01987_),
    .A2(_01836_),
    .B1(_01986_),
    .X(_02128_));
 sky130_fd_sc_hd__and2b_1 _21932_ (.A_N(_01992_),
    .B(_02014_),
    .X(_02129_));
 sky130_fd_sc_hd__and2b_1 _21933_ (.A_N(_01990_),
    .B(_02015_),
    .X(_02130_));
 sky130_fd_sc_hd__or2_1 _21934_ (.A(_14396_),
    .B(_01834_),
    .X(_02131_));
 sky130_fd_sc_hd__a21oi_4 _21935_ (.A1(_14567_),
    .A2(_02131_),
    .B1(_01987_),
    .Y(_02132_));
 sky130_fd_sc_hd__o21ba_1 _21936_ (.A1(_02129_),
    .A2(_02130_),
    .B1_N(_02132_),
    .X(_02133_));
 sky130_fd_sc_hd__or3b_1 _21937_ (.A(_02129_),
    .B(_02130_),
    .C_N(_02132_),
    .X(_02134_));
 sky130_fd_sc_hd__and2b_1 _21938_ (.A_N(_02133_),
    .B(_02134_),
    .X(_02135_));
 sky130_fd_sc_hd__buf_2 _21939_ (.A(_01994_),
    .X(_02136_));
 sky130_fd_sc_hd__buf_2 _21940_ (.A(_02136_),
    .X(_02137_));
 sky130_fd_sc_hd__nor2_1 _21941_ (.A(_02137_),
    .B(_02013_),
    .Y(_02138_));
 sky130_fd_sc_hd__a21o_1 _21942_ (.A1(_02011_),
    .A2(_02012_),
    .B1(_02138_),
    .X(_02139_));
 sky130_fd_sc_hd__or3b_1 _21943_ (.A(_02017_),
    .B(_02050_),
    .C_N(_02051_),
    .X(_02140_));
 sky130_fd_sc_hd__and2b_1 _21944_ (.A_N(_02050_),
    .B(_02140_),
    .X(_02141_));
 sky130_fd_sc_hd__or2b_1 _21945_ (.A(_02000_),
    .B_N(_02004_),
    .X(_02142_));
 sky130_fd_sc_hd__or2b_1 _21946_ (.A(_01999_),
    .B_N(_02005_),
    .X(_02143_));
 sky130_fd_sc_hd__a32o_2 _21947_ (.A1(_02028_),
    .A2(_02029_),
    .A3(_02031_),
    .B1(_02032_),
    .B2(_02024_),
    .X(_02144_));
 sky130_fd_sc_hd__o2bb2ai_1 _21948_ (.A1_N(_14212_),
    .A2_N(_02001_),
    .B1(_02003_),
    .B2(_01850_),
    .Y(_02145_));
 sky130_fd_sc_hd__and4_1 _21949_ (.A(_13661_),
    .B(_13662_),
    .C(_01516_),
    .D(_14033_),
    .X(_02146_));
 sky130_fd_sc_hd__o21ai_4 _21950_ (.A1(_10836_),
    .A2(_10839_),
    .B1(\genblk1.pcpi_mul.rs1[32] ),
    .Y(_02147_));
 sky130_fd_sc_hd__or3_1 _21951_ (.A(_01850_),
    .B(_02001_),
    .C(_02147_),
    .X(_02148_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _21952_ (.A(_02148_),
    .X(_02149_));
 sky130_fd_sc_hd__o21ai_1 _21953_ (.A1(_02001_),
    .A2(_02147_),
    .B1(_01850_),
    .Y(_02150_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _21954_ (.A(_02150_),
    .X(_02151_));
 sky130_fd_sc_hd__o211a_1 _21955_ (.A1(_02146_),
    .A2(_02023_),
    .B1(_02149_),
    .C1(_02151_),
    .X(_02152_));
 sky130_fd_sc_hd__a211oi_1 _21956_ (.A1(_02149_),
    .A2(_02151_),
    .B1(_02146_),
    .C1(_02023_),
    .Y(_02153_));
 sky130_fd_sc_hd__nor2_1 _21957_ (.A(_02152_),
    .B(_02153_),
    .Y(_02154_));
 sky130_fd_sc_hd__xor2_1 _21958_ (.A(_02145_),
    .B(_02154_),
    .X(_02155_));
 sky130_fd_sc_hd__xnor2_1 _21959_ (.A(_02144_),
    .B(_02155_),
    .Y(_02156_));
 sky130_fd_sc_hd__a21o_1 _21960_ (.A1(_02142_),
    .A2(_02143_),
    .B1(_02156_),
    .X(_02157_));
 sky130_fd_sc_hd__nand3_1 _21961_ (.A(_02142_),
    .B(_02143_),
    .C(_02156_),
    .Y(_02158_));
 sky130_fd_sc_hd__nand2_1 _21962_ (.A(_02157_),
    .B(_02158_),
    .Y(_02159_));
 sky130_fd_sc_hd__a21bo_1 _21963_ (.A1(_01997_),
    .A2(_02008_),
    .B1_N(_02007_),
    .X(_02160_));
 sky130_fd_sc_hd__xor2_1 _21964_ (.A(_02159_),
    .B(_02160_),
    .X(_02161_));
 sky130_fd_sc_hd__xor2_1 _21965_ (.A(_01995_),
    .B(_02161_),
    .X(_02162_));
 sky130_fd_sc_hd__xnor2_1 _21966_ (.A(_02141_),
    .B(_02162_),
    .Y(_02163_));
 sky130_fd_sc_hd__xnor2_1 _21967_ (.A(_02139_),
    .B(_02163_),
    .Y(_02164_));
 sky130_fd_sc_hd__nor2_2 _21968_ (.A(_02046_),
    .B(_02048_),
    .Y(_02165_));
 sky130_fd_sc_hd__a22oi_4 _21969_ (.A1(_11108_),
    .A2(_13608_),
    .B1(_13609_),
    .B2(_10957_),
    .Y(_02166_));
 sky130_fd_sc_hd__and4_1 _21970_ (.A(_10963_),
    .B(_11111_),
    .C(\genblk1.pcpi_mul.rs1[29] ),
    .D(\genblk1.pcpi_mul.rs1[30] ),
    .X(_02167_));
 sky130_fd_sc_hd__nor2_1 _21971_ (.A(_02166_),
    .B(_02167_),
    .Y(_02168_));
 sky130_fd_sc_hd__nand2_2 _21972_ (.A(_10961_),
    .B(_13618_),
    .Y(_02169_));
 sky130_fd_sc_hd__xnor2_2 _21973_ (.A(_02168_),
    .B(_02169_),
    .Y(_02170_));
 sky130_fd_sc_hd__a22oi_1 _21974_ (.A1(_14087_),
    .A2(_13867_),
    .B1(_13445_),
    .B2(_14086_),
    .Y(_02171_));
 sky130_fd_sc_hd__and4_1 _21975_ (.A(_11236_),
    .B(_13676_),
    .C(_12973_),
    .D(_12980_),
    .X(_02172_));
 sky130_fd_sc_hd__nor2_1 _21976_ (.A(_02171_),
    .B(_02172_),
    .Y(_02173_));
 sky130_fd_sc_hd__nand2_1 _21977_ (.A(_11135_),
    .B(_01516_),
    .Y(_02174_));
 sky130_fd_sc_hd__xnor2_2 _21978_ (.A(_02173_),
    .B(_02174_),
    .Y(_02175_));
 sky130_fd_sc_hd__nand2_1 _21979_ (.A(_02026_),
    .B(_02028_),
    .Y(_02176_));
 sky130_fd_sc_hd__xor2_1 _21980_ (.A(_02175_),
    .B(_02176_),
    .X(_02177_));
 sky130_fd_sc_hd__nand2_2 _21981_ (.A(_02170_),
    .B(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__or2_1 _21982_ (.A(_02170_),
    .B(_02177_),
    .X(_02179_));
 sky130_fd_sc_hd__nand2_1 _21983_ (.A(_02178_),
    .B(_02179_),
    .Y(_02180_));
 sky130_fd_sc_hd__or2b_1 _21984_ (.A(_02038_),
    .B_N(_02043_),
    .X(_02181_));
 sky130_fd_sc_hd__nand2_1 _21985_ (.A(_02037_),
    .B(_02044_),
    .Y(_02182_));
 sky130_fd_sc_hd__a31o_1 _21986_ (.A1(_11561_),
    .A2(_01544_),
    .A3(_02041_),
    .B1(_02040_),
    .X(_02183_));
 sky130_fd_sc_hd__o21ba_1 _21987_ (.A1(_02057_),
    .A2(_02059_),
    .B1_N(_02058_),
    .X(_02184_));
 sky130_fd_sc_hd__a22oi_1 _21988_ (.A1(_11781_),
    .A2(_12538_),
    .B1(_12690_),
    .B2(_11923_),
    .Y(_02185_));
 sky130_fd_sc_hd__and4_1 _21989_ (.A(_11662_),
    .B(_11658_),
    .C(_12537_),
    .D(_12688_),
    .X(_02186_));
 sky130_fd_sc_hd__nor2_1 _21990_ (.A(_02185_),
    .B(_02186_),
    .Y(_02187_));
 sky130_fd_sc_hd__nand2_1 _21991_ (.A(_11444_),
    .B(_13125_),
    .Y(_02188_));
 sky130_fd_sc_hd__xnor2_2 _21992_ (.A(_02187_),
    .B(_02188_),
    .Y(_02189_));
 sky130_fd_sc_hd__xnor2_1 _21993_ (.A(_02184_),
    .B(_02189_),
    .Y(_02190_));
 sky130_fd_sc_hd__xnor2_1 _21994_ (.A(_02183_),
    .B(_02190_),
    .Y(_02191_));
 sky130_fd_sc_hd__a21oi_1 _21995_ (.A1(_02181_),
    .A2(_02182_),
    .B1(_02191_),
    .Y(_02192_));
 sky130_fd_sc_hd__and3_1 _21996_ (.A(_02181_),
    .B(_02182_),
    .C(_02191_),
    .X(_02193_));
 sky130_fd_sc_hd__or3_1 _21997_ (.A(_02180_),
    .B(_02192_),
    .C(_02193_),
    .X(_02194_));
 sky130_fd_sc_hd__o21ai_1 _21998_ (.A1(_02192_),
    .A2(_02193_),
    .B1(_02180_),
    .Y(_02195_));
 sky130_fd_sc_hd__o211a_1 _21999_ (.A1(_02070_),
    .A2(_02072_),
    .B1(_02194_),
    .C1(_02195_),
    .X(_02196_));
 sky130_fd_sc_hd__a211o_1 _22000_ (.A1(_02194_),
    .A2(_02195_),
    .B1(_02070_),
    .C1(_02072_),
    .X(_02197_));
 sky130_fd_sc_hd__and2b_1 _22001_ (.A_N(_02196_),
    .B(_02197_),
    .X(_02198_));
 sky130_fd_sc_hd__xnor2_4 _22002_ (.A(_02165_),
    .B(_02198_),
    .Y(_02199_));
 sky130_fd_sc_hd__or2b_1 _22003_ (.A(_02067_),
    .B_N(_02066_),
    .X(_02200_));
 sky130_fd_sc_hd__nand2_1 _22004_ (.A(_02061_),
    .B(_02068_),
    .Y(_02201_));
 sky130_fd_sc_hd__or3_1 _22005_ (.A(_02075_),
    .B(_02078_),
    .C(_02079_),
    .X(_02202_));
 sky130_fd_sc_hd__a22oi_2 _22006_ (.A1(_01755_),
    .A2(_13663_),
    .B1(_12543_),
    .B2(_01754_),
    .Y(_02203_));
 sky130_fd_sc_hd__and4_1 _22007_ (.A(_14123_),
    .B(_12023_),
    .C(_13666_),
    .D(_14272_),
    .X(_02204_));
 sky130_fd_sc_hd__nor2_1 _22008_ (.A(_02203_),
    .B(_02204_),
    .Y(_02205_));
 sky130_fd_sc_hd__nand2_1 _22009_ (.A(_11771_),
    .B(_14269_),
    .Y(_02206_));
 sky130_fd_sc_hd__xnor2_2 _22010_ (.A(_02205_),
    .B(_02206_),
    .Y(_02207_));
 sky130_fd_sc_hd__a22oi_2 _22011_ (.A1(_11947_),
    .A2(_01912_),
    .B1(_13723_),
    .B2(_12074_),
    .Y(_02208_));
 sky130_fd_sc_hd__and4_1 _22012_ (.A(_12285_),
    .B(_11830_),
    .C(_14131_),
    .D(_13374_),
    .X(_02209_));
 sky130_fd_sc_hd__nor2_1 _22013_ (.A(_02208_),
    .B(_02209_),
    .Y(_02210_));
 sky130_fd_sc_hd__nand2_1 _22014_ (.A(_13674_),
    .B(_14482_),
    .Y(_02211_));
 sky130_fd_sc_hd__xnor2_1 _22015_ (.A(_02210_),
    .B(_02211_),
    .Y(_02212_));
 sky130_fd_sc_hd__o21ba_1 _22016_ (.A1(_02062_),
    .A2(_02064_),
    .B1_N(_02063_),
    .X(_02213_));
 sky130_fd_sc_hd__xnor2_1 _22017_ (.A(_02212_),
    .B(_02213_),
    .Y(_02214_));
 sky130_fd_sc_hd__xnor2_1 _22018_ (.A(_02207_),
    .B(_02214_),
    .Y(_02215_));
 sky130_fd_sc_hd__a21oi_1 _22019_ (.A1(_02202_),
    .A2(_02082_),
    .B1(_02215_),
    .Y(_02216_));
 sky130_fd_sc_hd__and3_1 _22020_ (.A(_02202_),
    .B(_02082_),
    .C(_02215_),
    .X(_02217_));
 sky130_fd_sc_hd__a211o_1 _22021_ (.A1(_02200_),
    .A2(_02201_),
    .B1(_02216_),
    .C1(_02217_),
    .X(_02218_));
 sky130_fd_sc_hd__o211ai_1 _22022_ (.A1(_02216_),
    .A2(_02217_),
    .B1(_02200_),
    .C1(_02201_),
    .Y(_02219_));
 sky130_fd_sc_hd__and2_2 _22023_ (.A(_02218_),
    .B(_02219_),
    .X(_02220_));
 sky130_fd_sc_hd__o21ba_1 _22024_ (.A1(_02085_),
    .A2(_02087_),
    .B1_N(_02086_),
    .X(_02221_));
 sky130_fd_sc_hd__a22oi_2 _22025_ (.A1(_11490_),
    .A2(_12771_),
    .B1(_13744_),
    .B2(_12561_),
    .Y(_02222_));
 sky130_fd_sc_hd__and4_2 _22026_ (.A(_11380_),
    .B(_11961_),
    .C(_13558_),
    .D(_13556_),
    .X(_02223_));
 sky130_fd_sc_hd__o2bb2a_1 _22027_ (.A1_N(_13690_),
    .A2_N(_12585_),
    .B1(_02222_),
    .B2(_02223_),
    .X(_02224_));
 sky130_fd_sc_hd__and4bb_1 _22028_ (.A_N(_02222_),
    .B_N(_02223_),
    .C(_13695_),
    .D(_14499_),
    .X(_02225_));
 sky130_fd_sc_hd__nor2_1 _22029_ (.A(_02224_),
    .B(_02225_),
    .Y(_02226_));
 sky130_fd_sc_hd__xnor2_1 _22030_ (.A(_02221_),
    .B(_02226_),
    .Y(_02227_));
 sky130_fd_sc_hd__o21ai_2 _22031_ (.A1(_02077_),
    .A2(_02079_),
    .B1(_02227_),
    .Y(_02228_));
 sky130_fd_sc_hd__or3_1 _22032_ (.A(_02077_),
    .B(_02079_),
    .C(_02227_),
    .X(_02229_));
 sky130_fd_sc_hd__and2_2 _22033_ (.A(_02228_),
    .B(_02229_),
    .X(_02230_));
 sky130_fd_sc_hd__nand2_1 _22034_ (.A(_11373_),
    .B(_14154_),
    .Y(_02231_));
 sky130_fd_sc_hd__and4_1 _22035_ (.A(_11160_),
    .B(_11261_),
    .C(_13760_),
    .D(_13971_),
    .X(_02232_));
 sky130_fd_sc_hd__a22oi_1 _22036_ (.A1(_11473_),
    .A2(_13228_),
    .B1(_13762_),
    .B2(_11728_),
    .Y(_02233_));
 sky130_fd_sc_hd__nor2_1 _22037_ (.A(_02232_),
    .B(_02233_),
    .Y(_02234_));
 sky130_fd_sc_hd__xnor2_2 _22038_ (.A(_02231_),
    .B(_02234_),
    .Y(_02235_));
 sky130_fd_sc_hd__nand2_1 _22039_ (.A(_11270_),
    .B(_14160_),
    .Y(_02236_));
 sky130_fd_sc_hd__buf_1 _22040_ (.A(\genblk1.pcpi_mul.rs2[32] ),
    .X(_02237_));
 sky130_fd_sc_hd__and2b_1 _22041_ (.A_N(_10858_),
    .B(_02237_),
    .X(_02238_));
 sky130_fd_sc_hd__nand2_1 _22042_ (.A(_11280_),
    .B(_14167_),
    .Y(_02239_));
 sky130_fd_sc_hd__xnor2_2 _22043_ (.A(_02238_),
    .B(_02239_),
    .Y(_02240_));
 sky130_fd_sc_hd__xnor2_2 _22044_ (.A(_02236_),
    .B(_02240_),
    .Y(_02241_));
 sky130_fd_sc_hd__and3_1 _22045_ (.A(_11049_),
    .B(_14168_),
    .C(_02091_),
    .X(_02242_));
 sky130_fd_sc_hd__a31o_1 _22046_ (.A1(_11167_),
    .A2(_14166_),
    .A3(_02093_),
    .B1(_02242_),
    .X(_02243_));
 sky130_fd_sc_hd__xor2_2 _22047_ (.A(_02241_),
    .B(_02243_),
    .X(_02244_));
 sky130_fd_sc_hd__xnor2_2 _22048_ (.A(_02235_),
    .B(_02244_),
    .Y(_02245_));
 sky130_fd_sc_hd__nand2_1 _22049_ (.A(_02094_),
    .B(_02096_),
    .Y(_02246_));
 sky130_fd_sc_hd__a21boi_4 _22050_ (.A1(_02089_),
    .A2(_02097_),
    .B1_N(_02246_),
    .Y(_02247_));
 sky130_fd_sc_hd__xnor2_2 _22051_ (.A(_02245_),
    .B(_02247_),
    .Y(_02248_));
 sky130_fd_sc_hd__xnor2_4 _22052_ (.A(_02230_),
    .B(_02248_),
    .Y(_02249_));
 sky130_fd_sc_hd__nand2_1 _22053_ (.A(_02098_),
    .B(_02100_),
    .Y(_02250_));
 sky130_fd_sc_hd__nor2_1 _22054_ (.A(_02098_),
    .B(_02100_),
    .Y(_02251_));
 sky130_fd_sc_hd__a21oi_4 _22055_ (.A1(_02084_),
    .A2(_02250_),
    .B1(_02251_),
    .Y(_02252_));
 sky130_fd_sc_hd__xnor2_4 _22056_ (.A(_02249_),
    .B(_02252_),
    .Y(_02253_));
 sky130_fd_sc_hd__xnor2_4 _22057_ (.A(_02220_),
    .B(_02253_),
    .Y(_02254_));
 sky130_fd_sc_hd__and2b_1 _22058_ (.A_N(_02105_),
    .B(_02102_),
    .X(_02255_));
 sky130_fd_sc_hd__a21oi_4 _22059_ (.A1(_02074_),
    .A2(_02106_),
    .B1(_02255_),
    .Y(_02256_));
 sky130_fd_sc_hd__xor2_4 _22060_ (.A(_02254_),
    .B(_02256_),
    .X(_02257_));
 sky130_fd_sc_hd__xor2_2 _22061_ (.A(_02199_),
    .B(_02257_),
    .X(_02258_));
 sky130_fd_sc_hd__nor2_1 _22062_ (.A(_02107_),
    .B(_02109_),
    .Y(_02259_));
 sky130_fd_sc_hd__a21o_1 _22063_ (.A1(_02053_),
    .A2(_02110_),
    .B1(_02259_),
    .X(_02260_));
 sky130_fd_sc_hd__xor2_1 _22064_ (.A(_02258_),
    .B(_02260_),
    .X(_02261_));
 sky130_fd_sc_hd__xnor2_1 _22065_ (.A(_02164_),
    .B(_02261_),
    .Y(_02262_));
 sky130_fd_sc_hd__and2b_1 _22066_ (.A_N(_02113_),
    .B(_02111_),
    .X(_02263_));
 sky130_fd_sc_hd__a21oi_1 _22067_ (.A1(_02016_),
    .A2(_02114_),
    .B1(_02263_),
    .Y(_02264_));
 sky130_fd_sc_hd__xnor2_1 _22068_ (.A(_02262_),
    .B(_02264_),
    .Y(_02265_));
 sky130_fd_sc_hd__xnor2_1 _22069_ (.A(_02135_),
    .B(_02265_),
    .Y(_02266_));
 sky130_fd_sc_hd__nor2_1 _22070_ (.A(_02115_),
    .B(_02117_),
    .Y(_02267_));
 sky130_fd_sc_hd__a21oi_1 _22071_ (.A1(_01989_),
    .A2(_02118_),
    .B1(_02267_),
    .Y(_02268_));
 sky130_fd_sc_hd__or2_1 _22072_ (.A(_02266_),
    .B(_02268_),
    .X(_02269_));
 sky130_fd_sc_hd__nand2_1 _22073_ (.A(_02266_),
    .B(_02268_),
    .Y(_02270_));
 sky130_fd_sc_hd__and2_1 _22074_ (.A(_02269_),
    .B(_02270_),
    .X(_02271_));
 sky130_fd_sc_hd__xnor2_1 _22075_ (.A(_02128_),
    .B(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hd__and2b_1 _22076_ (.A_N(_02121_),
    .B(_02119_),
    .X(_02273_));
 sky130_fd_sc_hd__a21oi_1 _22077_ (.A1(_01982_),
    .A2(_02122_),
    .B1(_02273_),
    .Y(_02274_));
 sky130_fd_sc_hd__nor2_1 _22078_ (.A(_02272_),
    .B(_02274_),
    .Y(_02275_));
 sky130_fd_sc_hd__and2_1 _22079_ (.A(_02272_),
    .B(_02274_),
    .X(_02276_));
 sky130_fd_sc_hd__or2_2 _22080_ (.A(_02275_),
    .B(_02276_),
    .X(_02277_));
 sky130_fd_sc_hd__and2_1 _22081_ (.A(_01976_),
    .B(_02124_),
    .X(_02278_));
 sky130_fd_sc_hd__a21o_1 _22082_ (.A1(_01981_),
    .A2(_02123_),
    .B1(_02125_),
    .X(_02279_));
 sky130_fd_sc_hd__o21ai_1 _22083_ (.A1(_01981_),
    .A2(_02123_),
    .B1(_02279_),
    .Y(_02280_));
 sky130_fd_sc_hd__a31o_1 _22084_ (.A1(_01824_),
    .A2(_01977_),
    .A3(_02278_),
    .B1(_02280_),
    .X(_02281_));
 sky130_fd_sc_hd__nand3b_2 _22085_ (.A_N(_01659_),
    .B(_01825_),
    .C(_02278_),
    .Y(_02282_));
 sky130_fd_sc_hd__nor2_2 _22086_ (.A(net334),
    .B(_02282_),
    .Y(_02283_));
 sky130_fd_sc_hd__a211oi_4 _22087_ (.A1(_14007_),
    .A2(_14009_),
    .B1(_01664_),
    .C1(_02282_),
    .Y(_02284_));
 sky130_fd_sc_hd__or3_2 _22088_ (.A(_02281_),
    .B(_02283_),
    .C(_02284_),
    .X(_02285_));
 sky130_fd_sc_hd__xnor2_4 _22089_ (.A(_02277_),
    .B(_02285_),
    .Y(_00086_));
 sky130_fd_sc_hd__nand2_1 _22090_ (.A(_02128_),
    .B(_02271_),
    .Y(_02286_));
 sky130_fd_sc_hd__buf_4 _22091_ (.A(_02132_),
    .X(_02287_));
 sky130_fd_sc_hd__and2b_1 _22092_ (.A_N(_02141_),
    .B(_02162_),
    .X(_02288_));
 sky130_fd_sc_hd__a21oi_2 _22093_ (.A1(_02139_),
    .A2(_02163_),
    .B1(_02288_),
    .Y(_02289_));
 sky130_fd_sc_hd__xnor2_2 _22094_ (.A(_02287_),
    .B(_02289_),
    .Y(_02290_));
 sky130_fd_sc_hd__nor2_1 _22095_ (.A(_02137_),
    .B(_02161_),
    .Y(_02291_));
 sky130_fd_sc_hd__a31o_1 _22096_ (.A1(_02157_),
    .A2(_02158_),
    .A3(_02160_),
    .B1(_02291_),
    .X(_02292_));
 sky130_fd_sc_hd__or3b_1 _22097_ (.A(_02165_),
    .B(_02196_),
    .C_N(_02197_),
    .X(_02293_));
 sky130_fd_sc_hd__or2b_1 _22098_ (.A(_02196_),
    .B_N(_02293_),
    .X(_02294_));
 sky130_fd_sc_hd__a21oi_2 _22099_ (.A1(_02145_),
    .A2(_02154_),
    .B1(_02152_),
    .Y(_02295_));
 sky130_fd_sc_hd__nand2_1 _22100_ (.A(_02175_),
    .B(_02176_),
    .Y(_02296_));
 sky130_fd_sc_hd__or2b_1 _22101_ (.A(_02001_),
    .B_N(_02148_),
    .X(_02297_));
 sky130_fd_sc_hd__clkbuf_2 _22102_ (.A(_02297_),
    .X(_02298_));
 sky130_fd_sc_hd__o21bai_4 _22103_ (.A1(_02166_),
    .A2(_02169_),
    .B1_N(_02167_),
    .Y(_02299_));
 sky130_fd_sc_hd__and3_1 _22104_ (.A(_02148_),
    .B(_02150_),
    .C(_02299_),
    .X(_02300_));
 sky130_fd_sc_hd__a21oi_1 _22105_ (.A1(_02149_),
    .A2(_02151_),
    .B1(_02299_),
    .Y(_02301_));
 sky130_fd_sc_hd__nor2_1 _22106_ (.A(_02300_),
    .B(_02301_),
    .Y(_02302_));
 sky130_fd_sc_hd__xnor2_1 _22107_ (.A(_02298_),
    .B(_02302_),
    .Y(_02303_));
 sky130_fd_sc_hd__a21oi_1 _22108_ (.A1(_02296_),
    .A2(_02178_),
    .B1(_02303_),
    .Y(_02304_));
 sky130_fd_sc_hd__and3_1 _22109_ (.A(_02296_),
    .B(_02178_),
    .C(_02303_),
    .X(_02305_));
 sky130_fd_sc_hd__or2_1 _22110_ (.A(_02304_),
    .B(_02305_),
    .X(_02306_));
 sky130_fd_sc_hd__xnor2_2 _22111_ (.A(_02295_),
    .B(_02306_),
    .Y(_02307_));
 sky130_fd_sc_hd__a21bo_1 _22112_ (.A1(_02144_),
    .A2(_02155_),
    .B1_N(_02157_),
    .X(_02308_));
 sky130_fd_sc_hd__xor2_2 _22113_ (.A(_02307_),
    .B(_02308_),
    .X(_02309_));
 sky130_fd_sc_hd__xor2_1 _22114_ (.A(_01995_),
    .B(_02309_),
    .X(_02310_));
 sky130_fd_sc_hd__xnor2_1 _22115_ (.A(_02294_),
    .B(_02310_),
    .Y(_02311_));
 sky130_fd_sc_hd__xnor2_2 _22116_ (.A(_02292_),
    .B(_02311_),
    .Y(_02312_));
 sky130_fd_sc_hd__and2b_2 _22117_ (.A_N(_02192_),
    .B(_02194_),
    .X(_02313_));
 sky130_fd_sc_hd__a21o_1 _22118_ (.A1(_02202_),
    .A2(_02082_),
    .B1(_02215_),
    .X(_02314_));
 sky130_fd_sc_hd__a22oi_2 _22119_ (.A1(_13662_),
    .A2(_14225_),
    .B1(_14210_),
    .B2(_13670_),
    .Y(_02315_));
 sky130_fd_sc_hd__and4_1 _22120_ (.A(_13661_),
    .B(_11112_),
    .C(_01846_),
    .D(_14398_),
    .X(_02316_));
 sky130_fd_sc_hd__or2_1 _22121_ (.A(_02315_),
    .B(_02316_),
    .X(_02317_));
 sky130_fd_sc_hd__nand2_4 _22122_ (.A(_11191_),
    .B(_14026_),
    .Y(_02318_));
 sky130_fd_sc_hd__xnor2_2 _22123_ (.A(_02317_),
    .B(_02318_),
    .Y(_02319_));
 sky130_fd_sc_hd__a22o_1 _22124_ (.A1(_13900_),
    .A2(_14417_),
    .B1(_14418_),
    .B2(_13680_),
    .X(_02320_));
 sky130_fd_sc_hd__nand4_2 _22125_ (.A(_11242_),
    .B(_13903_),
    .C(_13838_),
    .D(_13839_),
    .Y(_02321_));
 sky130_fd_sc_hd__a22o_1 _22126_ (.A1(_11233_),
    .A2(_13825_),
    .B1(_02320_),
    .B2(_02321_),
    .X(_02322_));
 sky130_fd_sc_hd__nand4_1 _22127_ (.A(_13897_),
    .B(_13814_),
    .C(_02320_),
    .D(_02321_),
    .Y(_02323_));
 sky130_fd_sc_hd__a31o_1 _22128_ (.A1(_11233_),
    .A2(_01717_),
    .A3(_02173_),
    .B1(_02172_),
    .X(_02324_));
 sky130_fd_sc_hd__and3_1 _22129_ (.A(_02322_),
    .B(_02323_),
    .C(_02324_),
    .X(_02325_));
 sky130_fd_sc_hd__a21oi_1 _22130_ (.A1(_02322_),
    .A2(_02323_),
    .B1(_02324_),
    .Y(_02326_));
 sky130_fd_sc_hd__nor2_1 _22131_ (.A(_02325_),
    .B(_02326_),
    .Y(_02327_));
 sky130_fd_sc_hd__xnor2_2 _22132_ (.A(_02319_),
    .B(_02327_),
    .Y(_02328_));
 sky130_fd_sc_hd__or2b_1 _22133_ (.A(_02184_),
    .B_N(_02189_),
    .X(_02329_));
 sky130_fd_sc_hd__nand2_1 _22134_ (.A(_02183_),
    .B(_02190_),
    .Y(_02330_));
 sky130_fd_sc_hd__buf_2 _22135_ (.A(_01540_),
    .X(_02331_));
 sky130_fd_sc_hd__a31o_1 _22136_ (.A1(_11446_),
    .A2(_02331_),
    .A3(_02187_),
    .B1(_02186_),
    .X(_02332_));
 sky130_fd_sc_hd__o21ba_1 _22137_ (.A1(_02203_),
    .A2(_02206_),
    .B1_N(_02204_),
    .X(_02333_));
 sky130_fd_sc_hd__a22oi_1 _22138_ (.A1(_11659_),
    .A2(_13859_),
    .B1(_13125_),
    .B2(_11656_),
    .Y(_02334_));
 sky130_fd_sc_hd__and4_1 _22139_ (.A(_11663_),
    .B(_13691_),
    .C(_12546_),
    .D(_13636_),
    .X(_02335_));
 sky130_fd_sc_hd__nor2_1 _22140_ (.A(_02334_),
    .B(_02335_),
    .Y(_02336_));
 sky130_fd_sc_hd__nand2_1 _22141_ (.A(_11775_),
    .B(_13286_),
    .Y(_02337_));
 sky130_fd_sc_hd__xnor2_2 _22142_ (.A(_02336_),
    .B(_02337_),
    .Y(_02338_));
 sky130_fd_sc_hd__xnor2_1 _22143_ (.A(_02333_),
    .B(_02338_),
    .Y(_02339_));
 sky130_fd_sc_hd__xnor2_1 _22144_ (.A(_02332_),
    .B(_02339_),
    .Y(_02340_));
 sky130_fd_sc_hd__a21o_1 _22145_ (.A1(_02329_),
    .A2(_02330_),
    .B1(_02340_),
    .X(_02341_));
 sky130_fd_sc_hd__nand3_1 _22146_ (.A(_02329_),
    .B(_02330_),
    .C(_02340_),
    .Y(_02342_));
 sky130_fd_sc_hd__and3_1 _22147_ (.A(_02328_),
    .B(_02341_),
    .C(_02342_),
    .X(_02343_));
 sky130_fd_sc_hd__a21oi_1 _22148_ (.A1(_02341_),
    .A2(_02342_),
    .B1(_02328_),
    .Y(_02344_));
 sky130_fd_sc_hd__a211oi_1 _22149_ (.A1(_02314_),
    .A2(_02218_),
    .B1(_02343_),
    .C1(_02344_),
    .Y(_02345_));
 sky130_fd_sc_hd__o211ai_1 _22150_ (.A1(_02343_),
    .A2(_02344_),
    .B1(_02314_),
    .C1(_02218_),
    .Y(_02346_));
 sky130_fd_sc_hd__and2b_1 _22151_ (.A_N(_02345_),
    .B(_02346_),
    .X(_02347_));
 sky130_fd_sc_hd__xnor2_4 _22152_ (.A(_02313_),
    .B(_02347_),
    .Y(_02348_));
 sky130_fd_sc_hd__or2b_1 _22153_ (.A(_02213_),
    .B_N(_02212_),
    .X(_02349_));
 sky130_fd_sc_hd__nand2_1 _22154_ (.A(_02207_),
    .B(_02214_),
    .Y(_02350_));
 sky130_fd_sc_hd__or3_1 _22155_ (.A(_02221_),
    .B(_02224_),
    .C(_02225_),
    .X(_02351_));
 sky130_fd_sc_hd__a22oi_2 _22156_ (.A1(_13716_),
    .A2(_12543_),
    .B1(_14269_),
    .B2(_01754_),
    .Y(_02352_));
 sky130_fd_sc_hd__and4_1 _22157_ (.A(_11896_),
    .B(_13934_),
    .C(_14272_),
    .D(_13890_),
    .X(_02353_));
 sky130_fd_sc_hd__nor2_1 _22158_ (.A(_02352_),
    .B(_02353_),
    .Y(_02354_));
 sky130_fd_sc_hd__nand2_1 _22159_ (.A(_11771_),
    .B(_14444_),
    .Y(_02355_));
 sky130_fd_sc_hd__xnor2_1 _22160_ (.A(_02354_),
    .B(_02355_),
    .Y(_02356_));
 sky130_fd_sc_hd__a22oi_2 _22161_ (.A1(_13305_),
    .A2(_01912_),
    .B1(_13723_),
    .B2(_11947_),
    .Y(_02357_));
 sky130_fd_sc_hd__and4_1 _22162_ (.A(_11830_),
    .B(_12067_),
    .C(_12328_),
    .D(_13374_),
    .X(_02358_));
 sky130_fd_sc_hd__nor2_1 _22163_ (.A(_02357_),
    .B(_02358_),
    .Y(_02359_));
 sky130_fd_sc_hd__nand2_1 _22164_ (.A(_13663_),
    .B(_14482_),
    .Y(_02360_));
 sky130_fd_sc_hd__xnor2_1 _22165_ (.A(_02359_),
    .B(_02360_),
    .Y(_02361_));
 sky130_fd_sc_hd__o21ba_1 _22166_ (.A1(_02208_),
    .A2(_02211_),
    .B1_N(_02209_),
    .X(_02362_));
 sky130_fd_sc_hd__xnor2_1 _22167_ (.A(_02361_),
    .B(_02362_),
    .Y(_02363_));
 sky130_fd_sc_hd__xnor2_1 _22168_ (.A(_02356_),
    .B(_02363_),
    .Y(_02364_));
 sky130_fd_sc_hd__a21oi_1 _22169_ (.A1(_02351_),
    .A2(_02228_),
    .B1(_02364_),
    .Y(_02365_));
 sky130_fd_sc_hd__and3_1 _22170_ (.A(_02351_),
    .B(_02228_),
    .C(_02364_),
    .X(_02366_));
 sky130_fd_sc_hd__a211o_1 _22171_ (.A1(_02349_),
    .A2(_02350_),
    .B1(_02365_),
    .C1(_02366_),
    .X(_02367_));
 sky130_fd_sc_hd__o211ai_1 _22172_ (.A1(_02365_),
    .A2(_02366_),
    .B1(_02349_),
    .C1(_02350_),
    .Y(_02368_));
 sky130_fd_sc_hd__and2_2 _22173_ (.A(_02367_),
    .B(_02368_),
    .X(_02369_));
 sky130_fd_sc_hd__o21ba_1 _22174_ (.A1(_02231_),
    .A2(_02233_),
    .B1_N(_02232_),
    .X(_02370_));
 sky130_fd_sc_hd__a22oi_2 _22175_ (.A1(_13689_),
    .A2(_12776_),
    .B1(_01601_),
    .B2(_11590_),
    .Y(_02371_));
 sky130_fd_sc_hd__and4_2 _22176_ (.A(_11489_),
    .B(_11698_),
    .C(_13060_),
    .D(_13061_),
    .X(_02372_));
 sky130_fd_sc_hd__o2bb2a_1 _22177_ (.A1_N(_13918_),
    .A2_N(_14499_),
    .B1(_02371_),
    .B2(_02372_),
    .X(_02373_));
 sky130_fd_sc_hd__and4bb_1 _22178_ (.A_N(_02371_),
    .B_N(_02372_),
    .C(_13918_),
    .D(_14324_),
    .X(_02374_));
 sky130_fd_sc_hd__nor2_1 _22179_ (.A(_02373_),
    .B(_02374_),
    .Y(_02375_));
 sky130_fd_sc_hd__xnor2_1 _22180_ (.A(_02370_),
    .B(_02375_),
    .Y(_02376_));
 sky130_fd_sc_hd__o21ai_2 _22181_ (.A1(_02223_),
    .A2(_02225_),
    .B1(_02376_),
    .Y(_02377_));
 sky130_fd_sc_hd__or3_1 _22182_ (.A(_02223_),
    .B(_02225_),
    .C(_02376_),
    .X(_02378_));
 sky130_fd_sc_hd__and2_2 _22183_ (.A(_02377_),
    .B(_02378_),
    .X(_02379_));
 sky130_fd_sc_hd__a22oi_2 _22184_ (.A1(_11479_),
    .A2(_13764_),
    .B1(_14508_),
    .B2(_11473_),
    .Y(_02380_));
 sky130_fd_sc_hd__and4_1 _22185_ (.A(_11261_),
    .B(_11277_),
    .C(_13760_),
    .D(_13545_),
    .X(_02381_));
 sky130_fd_sc_hd__nor2_1 _22186_ (.A(_02380_),
    .B(_02381_),
    .Y(_02382_));
 sky130_fd_sc_hd__nand2_1 _22187_ (.A(_11381_),
    .B(_14154_),
    .Y(_02383_));
 sky130_fd_sc_hd__xnor2_2 _22188_ (.A(_02382_),
    .B(_02383_),
    .Y(_02384_));
 sky130_fd_sc_hd__nand2_1 _22189_ (.A(_11056_),
    .B(_14342_),
    .Y(_02385_));
 sky130_fd_sc_hd__and2b_1 _22190_ (.A_N(_10919_),
    .B(_02237_),
    .X(_02386_));
 sky130_fd_sc_hd__nand2_1 _22191_ (.A(_11038_),
    .B(_14167_),
    .Y(_02387_));
 sky130_fd_sc_hd__xnor2_2 _22192_ (.A(_02386_),
    .B(_02387_),
    .Y(_02388_));
 sky130_fd_sc_hd__xnor2_2 _22193_ (.A(_02385_),
    .B(_02388_),
    .Y(_02389_));
 sky130_fd_sc_hd__and3_1 _22194_ (.A(_11042_),
    .B(_01620_),
    .C(_02238_),
    .X(_02390_));
 sky130_fd_sc_hd__a31o_1 _22195_ (.A1(_11157_),
    .A2(_14343_),
    .A3(_02240_),
    .B1(_02390_),
    .X(_02391_));
 sky130_fd_sc_hd__xor2_2 _22196_ (.A(_02389_),
    .B(_02391_),
    .X(_02392_));
 sky130_fd_sc_hd__xnor2_2 _22197_ (.A(_02384_),
    .B(_02392_),
    .Y(_02393_));
 sky130_fd_sc_hd__nand2_1 _22198_ (.A(_02241_),
    .B(_02243_),
    .Y(_02394_));
 sky130_fd_sc_hd__a21boi_2 _22199_ (.A1(_02235_),
    .A2(_02244_),
    .B1_N(_02394_),
    .Y(_02395_));
 sky130_fd_sc_hd__xnor2_2 _22200_ (.A(_02393_),
    .B(_02395_),
    .Y(_02396_));
 sky130_fd_sc_hd__xnor2_4 _22201_ (.A(_02379_),
    .B(_02396_),
    .Y(_02397_));
 sky130_fd_sc_hd__nand2_1 _22202_ (.A(_02245_),
    .B(_02247_),
    .Y(_02398_));
 sky130_fd_sc_hd__nor2_1 _22203_ (.A(_02245_),
    .B(_02247_),
    .Y(_02399_));
 sky130_fd_sc_hd__a21oi_4 _22204_ (.A1(_02230_),
    .A2(_02398_),
    .B1(_02399_),
    .Y(_02400_));
 sky130_fd_sc_hd__xnor2_4 _22205_ (.A(_02397_),
    .B(_02400_),
    .Y(_02401_));
 sky130_fd_sc_hd__xnor2_4 _22206_ (.A(_02369_),
    .B(_02401_),
    .Y(_02402_));
 sky130_fd_sc_hd__and2b_1 _22207_ (.A_N(_02252_),
    .B(_02249_),
    .X(_02403_));
 sky130_fd_sc_hd__a21oi_4 _22208_ (.A1(_02220_),
    .A2(_02253_),
    .B1(_02403_),
    .Y(_02404_));
 sky130_fd_sc_hd__xor2_4 _22209_ (.A(_02402_),
    .B(_02404_),
    .X(_02405_));
 sky130_fd_sc_hd__xnor2_4 _22210_ (.A(_02348_),
    .B(_02405_),
    .Y(_02406_));
 sky130_fd_sc_hd__nor2_1 _22211_ (.A(_02254_),
    .B(_02256_),
    .Y(_02407_));
 sky130_fd_sc_hd__a21oi_4 _22212_ (.A1(_02199_),
    .A2(_02257_),
    .B1(_02407_),
    .Y(_02408_));
 sky130_fd_sc_hd__xor2_2 _22213_ (.A(_02406_),
    .B(_02408_),
    .X(_02409_));
 sky130_fd_sc_hd__xnor2_2 _22214_ (.A(_02312_),
    .B(_02409_),
    .Y(_02410_));
 sky130_fd_sc_hd__nor2_1 _22215_ (.A(_02258_),
    .B(_02260_),
    .Y(_02411_));
 sky130_fd_sc_hd__nand2_1 _22216_ (.A(_02258_),
    .B(_02260_),
    .Y(_02412_));
 sky130_fd_sc_hd__o21a_1 _22217_ (.A1(_02164_),
    .A2(_02411_),
    .B1(_02412_),
    .X(_02413_));
 sky130_fd_sc_hd__xnor2_2 _22218_ (.A(_02410_),
    .B(_02413_),
    .Y(_02414_));
 sky130_fd_sc_hd__xor2_2 _22219_ (.A(_02290_),
    .B(_02414_),
    .X(_02415_));
 sky130_fd_sc_hd__and2b_1 _22220_ (.A_N(_02264_),
    .B(_02262_),
    .X(_02416_));
 sky130_fd_sc_hd__a21oi_2 _22221_ (.A1(_02135_),
    .A2(_02265_),
    .B1(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__xnor2_2 _22222_ (.A(_02415_),
    .B(_02417_),
    .Y(_02418_));
 sky130_fd_sc_hd__xnor2_1 _22223_ (.A(_02133_),
    .B(_02418_),
    .Y(_02419_));
 sky130_fd_sc_hd__a21oi_2 _22224_ (.A1(_02269_),
    .A2(_02286_),
    .B1(_02419_),
    .Y(_02420_));
 sky130_fd_sc_hd__and3_1 _22225_ (.A(_02269_),
    .B(_02286_),
    .C(_02419_),
    .X(_02421_));
 sky130_fd_sc_hd__nor2_2 _22226_ (.A(_02420_),
    .B(_02421_),
    .Y(_02422_));
 sky130_fd_sc_hd__and2b_1 _22227_ (.A_N(_02277_),
    .B(_02285_),
    .X(_02423_));
 sky130_fd_sc_hd__nor2_2 _22228_ (.A(_02275_),
    .B(_02423_),
    .Y(_02424_));
 sky130_fd_sc_hd__xnor2_4 _22229_ (.A(_02422_),
    .B(_02424_),
    .Y(_00087_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _22230_ (.A(_02132_),
    .X(_02425_));
 sky130_fd_sc_hd__clkbuf_2 _22231_ (.A(_02425_),
    .X(_02426_));
 sky130_fd_sc_hd__buf_4 _22232_ (.A(_02426_),
    .X(_02427_));
 sky130_fd_sc_hd__nor2_2 _22233_ (.A(_02427_),
    .B(_02289_),
    .Y(_02428_));
 sky130_fd_sc_hd__nand2_1 _22234_ (.A(_02294_),
    .B(_02310_),
    .Y(_02429_));
 sky130_fd_sc_hd__or2b_1 _22235_ (.A(_02311_),
    .B_N(_02292_),
    .X(_02430_));
 sky130_fd_sc_hd__nand2_1 _22236_ (.A(_02429_),
    .B(_02430_),
    .Y(_02431_));
 sky130_fd_sc_hd__xor2_2 _22237_ (.A(_02287_),
    .B(_02431_),
    .X(_02432_));
 sky130_fd_sc_hd__buf_2 _22238_ (.A(_01995_),
    .X(_02433_));
 sky130_fd_sc_hd__or2b_1 _22239_ (.A(_02307_),
    .B_N(_02308_),
    .X(_02434_));
 sky130_fd_sc_hd__o21ai_2 _22240_ (.A1(_02433_),
    .A2(_02309_),
    .B1(_02434_),
    .Y(_02435_));
 sky130_fd_sc_hd__or3b_1 _22241_ (.A(_02313_),
    .B(_02345_),
    .C_N(_02346_),
    .X(_02436_));
 sky130_fd_sc_hd__or2b_2 _22242_ (.A(_02345_),
    .B_N(_02436_),
    .X(_02437_));
 sky130_fd_sc_hd__o21bai_2 _22243_ (.A1(_02319_),
    .A2(_02326_),
    .B1_N(_02325_),
    .Y(_02438_));
 sky130_fd_sc_hd__and2_1 _22244_ (.A(_02148_),
    .B(_02150_),
    .X(_02439_));
 sky130_fd_sc_hd__clkbuf_2 _22245_ (.A(_02439_),
    .X(_02440_));
 sky130_fd_sc_hd__o21bai_2 _22246_ (.A1(_02315_),
    .A2(_02318_),
    .B1_N(_02316_),
    .Y(_02441_));
 sky130_fd_sc_hd__xor2_1 _22247_ (.A(_02440_),
    .B(_02441_),
    .X(_02442_));
 sky130_fd_sc_hd__xnor2_1 _22248_ (.A(_02298_),
    .B(_02442_),
    .Y(_02443_));
 sky130_fd_sc_hd__xnor2_1 _22249_ (.A(_02438_),
    .B(_02443_),
    .Y(_02444_));
 sky130_fd_sc_hd__clkbuf_2 _22250_ (.A(_02298_),
    .X(_02445_));
 sky130_fd_sc_hd__a21oi_1 _22251_ (.A1(_02445_),
    .A2(_02302_),
    .B1(_02300_),
    .Y(_02446_));
 sky130_fd_sc_hd__xor2_1 _22252_ (.A(_02444_),
    .B(_02446_),
    .X(_02447_));
 sky130_fd_sc_hd__a21o_1 _22253_ (.A1(_02296_),
    .A2(_02178_),
    .B1(_02303_),
    .X(_02448_));
 sky130_fd_sc_hd__o21a_1 _22254_ (.A1(_02295_),
    .A2(_02305_),
    .B1(_02448_),
    .X(_02449_));
 sky130_fd_sc_hd__nor2_1 _22255_ (.A(_02447_),
    .B(_02449_),
    .Y(_02450_));
 sky130_fd_sc_hd__and2_1 _22256_ (.A(_02447_),
    .B(_02449_),
    .X(_02451_));
 sky130_fd_sc_hd__nor2_1 _22257_ (.A(_02450_),
    .B(_02451_),
    .Y(_02452_));
 sky130_fd_sc_hd__xnor2_1 _22258_ (.A(_02136_),
    .B(_02452_),
    .Y(_02453_));
 sky130_fd_sc_hd__xnor2_1 _22259_ (.A(_02437_),
    .B(_02453_),
    .Y(_02454_));
 sky130_fd_sc_hd__xnor2_2 _22260_ (.A(_02435_),
    .B(_02454_),
    .Y(_02455_));
 sky130_fd_sc_hd__a21bo_2 _22261_ (.A1(_02328_),
    .A2(_02342_),
    .B1_N(_02341_),
    .X(_02456_));
 sky130_fd_sc_hd__a21o_1 _22262_ (.A1(_02351_),
    .A2(_02228_),
    .B1(_02364_),
    .X(_02457_));
 sky130_fd_sc_hd__and3_1 _22263_ (.A(_11142_),
    .B(_11145_),
    .C(\genblk1.pcpi_mul.rs1[32] ),
    .X(_02458_));
 sky130_fd_sc_hd__a22o_1 _22264_ (.A1(_11112_),
    .A2(_14398_),
    .B1(_13842_),
    .B2(_13669_),
    .X(_02459_));
 sky130_fd_sc_hd__a21bo_1 _22265_ (.A1(_13831_),
    .A2(_02458_),
    .B1_N(_02459_),
    .X(_02460_));
 sky130_fd_sc_hd__xor2_1 _22266_ (.A(_02318_),
    .B(_02460_),
    .X(_02461_));
 sky130_fd_sc_hd__a22oi_2 _22267_ (.A1(_13678_),
    .A2(_14418_),
    .B1(_13813_),
    .B2(_13680_),
    .Y(_02462_));
 sky130_fd_sc_hd__and4_1 _22268_ (.A(_11236_),
    .B(_13676_),
    .C(_13281_),
    .D(_13292_),
    .X(_02463_));
 sky130_fd_sc_hd__nor2_1 _22269_ (.A(_02462_),
    .B(_02463_),
    .Y(_02464_));
 sky130_fd_sc_hd__nand2_1 _22270_ (.A(_11136_),
    .B(_14225_),
    .Y(_02465_));
 sky130_fd_sc_hd__xnor2_1 _22271_ (.A(_02464_),
    .B(_02465_),
    .Y(_02466_));
 sky130_fd_sc_hd__nand2_1 _22272_ (.A(_02321_),
    .B(_02323_),
    .Y(_02467_));
 sky130_fd_sc_hd__xor2_1 _22273_ (.A(_02466_),
    .B(_02467_),
    .X(_02468_));
 sky130_fd_sc_hd__xnor2_1 _22274_ (.A(_02461_),
    .B(_02468_),
    .Y(_02469_));
 sky130_fd_sc_hd__or2b_1 _22275_ (.A(_02333_),
    .B_N(_02338_),
    .X(_02470_));
 sky130_fd_sc_hd__nand2_1 _22276_ (.A(_02332_),
    .B(_02339_),
    .Y(_02471_));
 sky130_fd_sc_hd__buf_2 _22277_ (.A(_01538_),
    .X(_02472_));
 sky130_fd_sc_hd__a31o_1 _22278_ (.A1(_14099_),
    .A2(_02472_),
    .A3(_02336_),
    .B1(_02335_),
    .X(_02473_));
 sky130_fd_sc_hd__o21ba_1 _22279_ (.A1(_02352_),
    .A2(_02355_),
    .B1_N(_02353_),
    .X(_02474_));
 sky130_fd_sc_hd__a22oi_1 _22280_ (.A1(_11659_),
    .A2(_13632_),
    .B1(_13285_),
    .B2(_11656_),
    .Y(_02475_));
 sky130_fd_sc_hd__and4_1 _22281_ (.A(_14103_),
    .B(_13691_),
    .C(_13636_),
    .D(_13867_),
    .X(_02476_));
 sky130_fd_sc_hd__nor2_1 _22282_ (.A(_02475_),
    .B(_02476_),
    .Y(_02477_));
 sky130_fd_sc_hd__nand2_1 _22283_ (.A(_11775_),
    .B(_01713_),
    .Y(_02478_));
 sky130_fd_sc_hd__xnor2_1 _22284_ (.A(_02477_),
    .B(_02478_),
    .Y(_02479_));
 sky130_fd_sc_hd__xnor2_1 _22285_ (.A(_02474_),
    .B(_02479_),
    .Y(_02480_));
 sky130_fd_sc_hd__xnor2_1 _22286_ (.A(_02473_),
    .B(_02480_),
    .Y(_02481_));
 sky130_fd_sc_hd__a21oi_2 _22287_ (.A1(_02470_),
    .A2(_02471_),
    .B1(_02481_),
    .Y(_02482_));
 sky130_fd_sc_hd__and3_1 _22288_ (.A(_02470_),
    .B(_02471_),
    .C(_02481_),
    .X(_02483_));
 sky130_fd_sc_hd__nor3_1 _22289_ (.A(_02469_),
    .B(_02482_),
    .C(_02483_),
    .Y(_02484_));
 sky130_fd_sc_hd__o21a_1 _22290_ (.A1(_02482_),
    .A2(_02483_),
    .B1(_02469_),
    .X(_02485_));
 sky130_fd_sc_hd__a211oi_1 _22291_ (.A1(_02457_),
    .A2(_02367_),
    .B1(net359),
    .C1(_02485_),
    .Y(_02486_));
 sky130_fd_sc_hd__o211ai_2 _22292_ (.A1(net359),
    .A2(_02485_),
    .B1(_02457_),
    .C1(_02367_),
    .Y(_02487_));
 sky130_fd_sc_hd__or2b_1 _22293_ (.A(_02486_),
    .B_N(_02487_),
    .X(_02488_));
 sky130_fd_sc_hd__xnor2_2 _22294_ (.A(_02456_),
    .B(_02488_),
    .Y(_02489_));
 sky130_fd_sc_hd__or2b_1 _22295_ (.A(_02362_),
    .B_N(_02361_),
    .X(_02490_));
 sky130_fd_sc_hd__nand2_1 _22296_ (.A(_02356_),
    .B(_02363_),
    .Y(_02491_));
 sky130_fd_sc_hd__or3_1 _22297_ (.A(_02370_),
    .B(_02373_),
    .C(_02374_),
    .X(_02492_));
 sky130_fd_sc_hd__a22oi_2 _22298_ (.A1(_13716_),
    .A2(_13890_),
    .B1(_13887_),
    .B2(_11891_),
    .Y(_02493_));
 sky130_fd_sc_hd__and4_1 _22299_ (.A(_14123_),
    .B(_12023_),
    .C(_14268_),
    .D(_12830_),
    .X(_02494_));
 sky130_fd_sc_hd__nor2_1 _22300_ (.A(_02493_),
    .B(_02494_),
    .Y(_02495_));
 sky130_fd_sc_hd__nand2_1 _22301_ (.A(_11771_),
    .B(_13860_),
    .Y(_02496_));
 sky130_fd_sc_hd__xnor2_1 _22302_ (.A(_02495_),
    .B(_02496_),
    .Y(_02497_));
 sky130_fd_sc_hd__a22oi_2 _22303_ (.A1(_12147_),
    .A2(_14131_),
    .B1(_13944_),
    .B2(_13305_),
    .Y(_02498_));
 sky130_fd_sc_hd__and4_1 _22304_ (.A(_12067_),
    .B(_12144_),
    .C(_12328_),
    .D(_13376_),
    .X(_02499_));
 sky130_fd_sc_hd__nor2_1 _22305_ (.A(_02498_),
    .B(_02499_),
    .Y(_02500_));
 sky130_fd_sc_hd__nand2_1 _22306_ (.A(_14482_),
    .B(_14272_),
    .Y(_02501_));
 sky130_fd_sc_hd__xnor2_1 _22307_ (.A(_02500_),
    .B(_02501_),
    .Y(_02502_));
 sky130_fd_sc_hd__o21ba_1 _22308_ (.A1(_02357_),
    .A2(_02360_),
    .B1_N(_02358_),
    .X(_02503_));
 sky130_fd_sc_hd__xnor2_1 _22309_ (.A(_02502_),
    .B(_02503_),
    .Y(_02504_));
 sky130_fd_sc_hd__xnor2_1 _22310_ (.A(_02497_),
    .B(_02504_),
    .Y(_02505_));
 sky130_fd_sc_hd__a21oi_1 _22311_ (.A1(_02492_),
    .A2(_02377_),
    .B1(_02505_),
    .Y(_02506_));
 sky130_fd_sc_hd__and3_1 _22312_ (.A(_02492_),
    .B(_02377_),
    .C(_02505_),
    .X(_02507_));
 sky130_fd_sc_hd__a211o_1 _22313_ (.A1(_02490_),
    .A2(_02491_),
    .B1(_02506_),
    .C1(_02507_),
    .X(_02508_));
 sky130_fd_sc_hd__o211ai_1 _22314_ (.A1(_02506_),
    .A2(_02507_),
    .B1(_02490_),
    .C1(_02491_),
    .Y(_02509_));
 sky130_fd_sc_hd__and2_2 _22315_ (.A(_02508_),
    .B(_02509_),
    .X(_02510_));
 sky130_fd_sc_hd__o21ba_1 _22316_ (.A1(_02380_),
    .A2(_02383_),
    .B1_N(_02381_),
    .X(_02511_));
 sky130_fd_sc_hd__a22oi_2 _22317_ (.A1(_11819_),
    .A2(_13555_),
    .B1(_01601_),
    .B2(_11598_),
    .Y(_02512_));
 sky130_fd_sc_hd__and4_2 _22318_ (.A(_11698_),
    .B(_11707_),
    .C(_13060_),
    .D(_13061_),
    .X(_02513_));
 sky130_fd_sc_hd__o2bb2a_1 _22319_ (.A1_N(_11831_),
    .A2_N(_14324_),
    .B1(_02512_),
    .B2(_02513_),
    .X(_02514_));
 sky130_fd_sc_hd__and4bb_1 _22320_ (.A_N(_02512_),
    .B_N(_02513_),
    .C(_13679_),
    .D(_12584_),
    .X(_02515_));
 sky130_fd_sc_hd__nor2_1 _22321_ (.A(_02514_),
    .B(_02515_),
    .Y(_02516_));
 sky130_fd_sc_hd__xnor2_1 _22322_ (.A(_02511_),
    .B(_02516_),
    .Y(_02517_));
 sky130_fd_sc_hd__o21ai_2 _22323_ (.A1(_02372_),
    .A2(_02374_),
    .B1(_02517_),
    .Y(_02518_));
 sky130_fd_sc_hd__or3_1 _22324_ (.A(_02372_),
    .B(_02374_),
    .C(_02517_),
    .X(_02519_));
 sky130_fd_sc_hd__and2_2 _22325_ (.A(_02518_),
    .B(_02519_),
    .X(_02520_));
 sky130_fd_sc_hd__a22oi_1 _22326_ (.A1(_11381_),
    .A2(_13228_),
    .B1(_13762_),
    .B2(_11373_),
    .Y(_02521_));
 sky130_fd_sc_hd__and4_1 _22327_ (.A(_12343_),
    .B(_11834_),
    .C(_13223_),
    .D(_13971_),
    .X(_02522_));
 sky130_fd_sc_hd__nor2_1 _22328_ (.A(_02521_),
    .B(_02522_),
    .Y(_02523_));
 sky130_fd_sc_hd__nand2_1 _22329_ (.A(_11591_),
    .B(_14154_),
    .Y(_02524_));
 sky130_fd_sc_hd__xnor2_2 _22330_ (.A(_02523_),
    .B(_02524_),
    .Y(_02525_));
 sky130_fd_sc_hd__nand2_1 _22331_ (.A(_11473_),
    .B(_14342_),
    .Y(_02526_));
 sky130_fd_sc_hd__and2b_1 _22332_ (.A_N(_11268_),
    .B(_02237_),
    .X(_02527_));
 sky130_fd_sc_hd__nand2_1 _22333_ (.A(_11067_),
    .B(\genblk1.pcpi_mul.rs2[31] ),
    .Y(_02528_));
 sky130_fd_sc_hd__xnor2_2 _22334_ (.A(_02527_),
    .B(_02528_),
    .Y(_02529_));
 sky130_fd_sc_hd__xnor2_2 _22335_ (.A(_02526_),
    .B(_02529_),
    .Y(_02530_));
 sky130_fd_sc_hd__and3_1 _22336_ (.A(_11156_),
    .B(_13753_),
    .C(_02386_),
    .X(_02531_));
 sky130_fd_sc_hd__a31o_1 _22337_ (.A1(_11068_),
    .A2(_14160_),
    .A3(_02388_),
    .B1(_02531_),
    .X(_02532_));
 sky130_fd_sc_hd__xor2_2 _22338_ (.A(_02530_),
    .B(_02532_),
    .X(_02533_));
 sky130_fd_sc_hd__xnor2_2 _22339_ (.A(_02525_),
    .B(_02533_),
    .Y(_02534_));
 sky130_fd_sc_hd__nand2_1 _22340_ (.A(_02389_),
    .B(_02391_),
    .Y(_02535_));
 sky130_fd_sc_hd__a21boi_2 _22341_ (.A1(_02384_),
    .A2(_02392_),
    .B1_N(_02535_),
    .Y(_02536_));
 sky130_fd_sc_hd__xnor2_2 _22342_ (.A(_02534_),
    .B(_02536_),
    .Y(_02537_));
 sky130_fd_sc_hd__xnor2_4 _22343_ (.A(_02520_),
    .B(_02537_),
    .Y(_02538_));
 sky130_fd_sc_hd__nand2_1 _22344_ (.A(_02393_),
    .B(_02395_),
    .Y(_02539_));
 sky130_fd_sc_hd__nor2_1 _22345_ (.A(_02393_),
    .B(_02395_),
    .Y(_02540_));
 sky130_fd_sc_hd__a21oi_4 _22346_ (.A1(_02379_),
    .A2(_02539_),
    .B1(_02540_),
    .Y(_02541_));
 sky130_fd_sc_hd__xnor2_4 _22347_ (.A(_02538_),
    .B(_02541_),
    .Y(_02542_));
 sky130_fd_sc_hd__xnor2_4 _22348_ (.A(_02510_),
    .B(_02542_),
    .Y(_02543_));
 sky130_fd_sc_hd__and2b_1 _22349_ (.A_N(_02400_),
    .B(_02397_),
    .X(_02544_));
 sky130_fd_sc_hd__a21oi_2 _22350_ (.A1(_02369_),
    .A2(_02401_),
    .B1(_02544_),
    .Y(_02545_));
 sky130_fd_sc_hd__xor2_2 _22351_ (.A(_02543_),
    .B(_02545_),
    .X(_02546_));
 sky130_fd_sc_hd__xor2_2 _22352_ (.A(_02489_),
    .B(_02546_),
    .X(_02547_));
 sky130_fd_sc_hd__nor2_1 _22353_ (.A(_02402_),
    .B(_02404_),
    .Y(_02548_));
 sky130_fd_sc_hd__a21oi_2 _22354_ (.A1(_02348_),
    .A2(_02405_),
    .B1(_02548_),
    .Y(_02549_));
 sky130_fd_sc_hd__xnor2_2 _22355_ (.A(_02547_),
    .B(_02549_),
    .Y(_02550_));
 sky130_fd_sc_hd__xor2_2 _22356_ (.A(_02455_),
    .B(_02550_),
    .X(_02551_));
 sky130_fd_sc_hd__nor2_1 _22357_ (.A(_02406_),
    .B(_02408_),
    .Y(_02552_));
 sky130_fd_sc_hd__a21o_1 _22358_ (.A1(_02312_),
    .A2(_02409_),
    .B1(_02552_),
    .X(_02553_));
 sky130_fd_sc_hd__xor2_1 _22359_ (.A(_02551_),
    .B(_02553_),
    .X(_02554_));
 sky130_fd_sc_hd__xnor2_2 _22360_ (.A(_02432_),
    .B(_02554_),
    .Y(_02555_));
 sky130_fd_sc_hd__or2_1 _22361_ (.A(_02410_),
    .B(_02413_),
    .X(_02556_));
 sky130_fd_sc_hd__o21a_2 _22362_ (.A1(_02290_),
    .A2(_02414_),
    .B1(_02556_),
    .X(_02557_));
 sky130_fd_sc_hd__xnor2_4 _22363_ (.A(_02555_),
    .B(_02557_),
    .Y(_02558_));
 sky130_fd_sc_hd__xnor2_4 _22364_ (.A(_02428_),
    .B(_02558_),
    .Y(_02559_));
 sky130_fd_sc_hd__or2b_1 _22365_ (.A(_02417_),
    .B_N(_02415_),
    .X(_02560_));
 sky130_fd_sc_hd__a21boi_4 _22366_ (.A1(_02133_),
    .A2(_02418_),
    .B1_N(_02560_),
    .Y(_02561_));
 sky130_fd_sc_hd__xor2_4 _22367_ (.A(_02559_),
    .B(_02561_),
    .X(_02562_));
 sky130_fd_sc_hd__o21bai_2 _22368_ (.A1(_02275_),
    .A2(_02420_),
    .B1_N(_02421_),
    .Y(_02563_));
 sky130_fd_sc_hd__a21bo_4 _22369_ (.A1(_02423_),
    .A2(_02422_),
    .B1_N(_02563_),
    .X(_02564_));
 sky130_fd_sc_hd__xor2_4 _22370_ (.A(_02562_),
    .B(_02564_),
    .X(_00088_));
 sky130_fd_sc_hd__or2b_1 _22371_ (.A(_02557_),
    .B_N(_02555_),
    .X(_02565_));
 sky130_fd_sc_hd__a21boi_4 _22372_ (.A1(_02428_),
    .A2(_02558_),
    .B1_N(_02565_),
    .Y(_02566_));
 sky130_fd_sc_hd__clkbuf_4 _22373_ (.A(_02426_),
    .X(_02567_));
 sky130_fd_sc_hd__a21oi_4 _22374_ (.A1(_02429_),
    .A2(_02430_),
    .B1(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__nand2_1 _22375_ (.A(_02437_),
    .B(_02453_),
    .Y(_02569_));
 sky130_fd_sc_hd__or2b_1 _22376_ (.A(_02454_),
    .B_N(_02435_),
    .X(_02570_));
 sky130_fd_sc_hd__nand2_2 _22377_ (.A(_02569_),
    .B(_02570_),
    .Y(_02571_));
 sky130_fd_sc_hd__xnor2_4 _22378_ (.A(_02287_),
    .B(_02571_),
    .Y(_02572_));
 sky130_fd_sc_hd__o21ba_2 _22379_ (.A1(_02433_),
    .A2(_02451_),
    .B1_N(_02450_),
    .X(_02573_));
 sky130_fd_sc_hd__a21oi_2 _22380_ (.A1(_02456_),
    .A2(_02487_),
    .B1(_02486_),
    .Y(_02574_));
 sky130_fd_sc_hd__and2_1 _22381_ (.A(_02466_),
    .B(_02467_),
    .X(_02575_));
 sky130_fd_sc_hd__a21o_1 _22382_ (.A1(_02461_),
    .A2(_02468_),
    .B1(_02575_),
    .X(_02576_));
 sky130_fd_sc_hd__a32o_1 _22383_ (.A1(_10894_),
    .A2(_14037_),
    .A3(_02459_),
    .B1(_02458_),
    .B2(_13831_),
    .X(_02577_));
 sky130_fd_sc_hd__xor2_1 _22384_ (.A(_02440_),
    .B(_02577_),
    .X(_02578_));
 sky130_fd_sc_hd__xnor2_1 _22385_ (.A(_02298_),
    .B(_02578_),
    .Y(_02579_));
 sky130_fd_sc_hd__xor2_1 _22386_ (.A(_02576_),
    .B(_02579_),
    .X(_02580_));
 sky130_fd_sc_hd__and3_1 _22387_ (.A(_02149_),
    .B(_02151_),
    .C(_02441_),
    .X(_02581_));
 sky130_fd_sc_hd__a21oi_1 _22388_ (.A1(_02445_),
    .A2(_02442_),
    .B1(_02581_),
    .Y(_02582_));
 sky130_fd_sc_hd__or2_1 _22389_ (.A(_02580_),
    .B(_02582_),
    .X(_02583_));
 sky130_fd_sc_hd__nand2_1 _22390_ (.A(_02580_),
    .B(_02582_),
    .Y(_02584_));
 sky130_fd_sc_hd__and2_1 _22391_ (.A(_02583_),
    .B(_02584_),
    .X(_02585_));
 sky130_fd_sc_hd__and2b_1 _22392_ (.A_N(_02443_),
    .B(_02438_),
    .X(_02586_));
 sky130_fd_sc_hd__and2b_1 _22393_ (.A_N(_02446_),
    .B(_02444_),
    .X(_02587_));
 sky130_fd_sc_hd__nor2_1 _22394_ (.A(_02586_),
    .B(_02587_),
    .Y(_02588_));
 sky130_fd_sc_hd__xor2_2 _22395_ (.A(_02585_),
    .B(_02588_),
    .X(_02589_));
 sky130_fd_sc_hd__xor2_2 _22396_ (.A(_01995_),
    .B(_02589_),
    .X(_02590_));
 sky130_fd_sc_hd__xnor2_2 _22397_ (.A(_02574_),
    .B(_02590_),
    .Y(_02591_));
 sky130_fd_sc_hd__xnor2_4 _22398_ (.A(_02573_),
    .B(_02591_),
    .Y(_02592_));
 sky130_fd_sc_hd__nor2_2 _22399_ (.A(_02482_),
    .B(_02484_),
    .Y(_02593_));
 sky130_fd_sc_hd__a21o_1 _22400_ (.A1(_02492_),
    .A2(_02377_),
    .B1(_02505_),
    .X(_02594_));
 sky130_fd_sc_hd__or2_1 _22401_ (.A(_11142_),
    .B(_11111_),
    .X(_02595_));
 sky130_fd_sc_hd__and3b_1 _22402_ (.A_N(_02458_),
    .B(_02595_),
    .C(_14570_),
    .X(_02596_));
 sky130_fd_sc_hd__xnor2_2 _22403_ (.A(_02318_),
    .B(_02596_),
    .Y(_02597_));
 sky130_fd_sc_hd__buf_4 _22404_ (.A(_02597_),
    .X(_02598_));
 sky130_fd_sc_hd__a22oi_1 _22405_ (.A1(_13903_),
    .A2(_13813_),
    .B1(_01846_),
    .B2(_11242_),
    .Y(_02599_));
 sky130_fd_sc_hd__and4_1 _22406_ (.A(_13680_),
    .B(_13678_),
    .C(_13608_),
    .D(_13609_),
    .X(_02600_));
 sky130_fd_sc_hd__o2bb2a_1 _22407_ (.A1_N(_13897_),
    .A2_N(_13827_),
    .B1(_02599_),
    .B2(_02600_),
    .X(_02601_));
 sky130_fd_sc_hd__and4bb_1 _22408_ (.A_N(_02599_),
    .B_N(_02600_),
    .C(_13897_),
    .D(_14210_),
    .X(_02602_));
 sky130_fd_sc_hd__o21ba_1 _22409_ (.A1(_02462_),
    .A2(_02465_),
    .B1_N(_02463_),
    .X(_02603_));
 sky130_fd_sc_hd__or3_1 _22410_ (.A(_02601_),
    .B(_02602_),
    .C(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__o21ai_1 _22411_ (.A1(_02601_),
    .A2(_02602_),
    .B1(_02603_),
    .Y(_02605_));
 sky130_fd_sc_hd__and2_1 _22412_ (.A(_02604_),
    .B(_02605_),
    .X(_02606_));
 sky130_fd_sc_hd__xnor2_1 _22413_ (.A(_02598_),
    .B(_02606_),
    .Y(_02607_));
 sky130_fd_sc_hd__or2b_1 _22414_ (.A(_02474_),
    .B_N(_02479_),
    .X(_02608_));
 sky130_fd_sc_hd__nand2_1 _22415_ (.A(_02473_),
    .B(_02480_),
    .Y(_02609_));
 sky130_fd_sc_hd__buf_2 _22416_ (.A(_01713_),
    .X(_02610_));
 sky130_fd_sc_hd__a31o_2 _22417_ (.A1(_11446_),
    .A2(_02610_),
    .A3(_02477_),
    .B1(_02476_),
    .X(_02611_));
 sky130_fd_sc_hd__o21ba_1 _22418_ (.A1(_02493_),
    .A2(_02496_),
    .B1_N(_02494_),
    .X(_02612_));
 sky130_fd_sc_hd__a22oi_2 _22419_ (.A1(_11659_),
    .A2(_13867_),
    .B1(_14417_),
    .B2(_11556_),
    .Y(_02613_));
 sky130_fd_sc_hd__and4_1 _22420_ (.A(_11663_),
    .B(_11925_),
    .C(_13867_),
    .D(_13445_),
    .X(_02614_));
 sky130_fd_sc_hd__nor2_1 _22421_ (.A(_02613_),
    .B(_02614_),
    .Y(_02615_));
 sky130_fd_sc_hd__nand2_1 _22422_ (.A(_11560_),
    .B(_13836_),
    .Y(_02616_));
 sky130_fd_sc_hd__xnor2_2 _22423_ (.A(_02615_),
    .B(_02616_),
    .Y(_02617_));
 sky130_fd_sc_hd__xnor2_1 _22424_ (.A(_02612_),
    .B(_02617_),
    .Y(_02618_));
 sky130_fd_sc_hd__xnor2_1 _22425_ (.A(_02611_),
    .B(_02618_),
    .Y(_02619_));
 sky130_fd_sc_hd__a21oi_1 _22426_ (.A1(_02608_),
    .A2(_02609_),
    .B1(_02619_),
    .Y(_02620_));
 sky130_fd_sc_hd__and3_1 _22427_ (.A(_02608_),
    .B(_02609_),
    .C(_02619_),
    .X(_02621_));
 sky130_fd_sc_hd__nor3_1 _22428_ (.A(_02607_),
    .B(_02620_),
    .C(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__o21a_1 _22429_ (.A1(_02620_),
    .A2(_02621_),
    .B1(_02607_),
    .X(_02623_));
 sky130_fd_sc_hd__a211oi_1 _22430_ (.A1(_02594_),
    .A2(_02508_),
    .B1(_02622_),
    .C1(_02623_),
    .Y(_02624_));
 sky130_fd_sc_hd__o211ai_1 _22431_ (.A1(_02622_),
    .A2(_02623_),
    .B1(_02594_),
    .C1(_02508_),
    .Y(_02625_));
 sky130_fd_sc_hd__and2b_1 _22432_ (.A_N(_02624_),
    .B(_02625_),
    .X(_02626_));
 sky130_fd_sc_hd__xnor2_4 _22433_ (.A(_02593_),
    .B(_02626_),
    .Y(_02627_));
 sky130_fd_sc_hd__or2b_1 _22434_ (.A(_02503_),
    .B_N(_02502_),
    .X(_02628_));
 sky130_fd_sc_hd__nand2_1 _22435_ (.A(_02497_),
    .B(_02504_),
    .Y(_02629_));
 sky130_fd_sc_hd__or3_1 _22436_ (.A(_02511_),
    .B(_02514_),
    .C(_02515_),
    .X(_02630_));
 sky130_fd_sc_hd__a22oi_1 _22437_ (.A1(_01755_),
    .A2(_14444_),
    .B1(_13860_),
    .B2(_01754_),
    .Y(_02631_));
 sky130_fd_sc_hd__and4_1 _22438_ (.A(_11896_),
    .B(_13934_),
    .C(_14080_),
    .D(_14076_),
    .X(_02632_));
 sky130_fd_sc_hd__nor2_1 _22439_ (.A(_02631_),
    .B(_02632_),
    .Y(_02633_));
 sky130_fd_sc_hd__nand2_1 _22440_ (.A(_13711_),
    .B(_13861_),
    .Y(_02634_));
 sky130_fd_sc_hd__xnor2_1 _22441_ (.A(_02633_),
    .B(_02634_),
    .Y(_02635_));
 sky130_fd_sc_hd__a22oi_2 _22442_ (.A1(_12154_),
    .A2(_01912_),
    .B1(_13723_),
    .B2(_12079_),
    .Y(_02636_));
 sky130_fd_sc_hd__and4_1 _22443_ (.A(_12147_),
    .B(_12271_),
    .C(_14131_),
    .D(_13374_),
    .X(_02637_));
 sky130_fd_sc_hd__nor2_1 _22444_ (.A(_02636_),
    .B(_02637_),
    .Y(_02638_));
 sky130_fd_sc_hd__nand2_1 _22445_ (.A(_14482_),
    .B(_13890_),
    .Y(_02639_));
 sky130_fd_sc_hd__xnor2_1 _22446_ (.A(_02638_),
    .B(_02639_),
    .Y(_02640_));
 sky130_fd_sc_hd__o21ba_1 _22447_ (.A1(_02498_),
    .A2(_02501_),
    .B1_N(_02499_),
    .X(_02641_));
 sky130_fd_sc_hd__xnor2_1 _22448_ (.A(_02640_),
    .B(_02641_),
    .Y(_02642_));
 sky130_fd_sc_hd__xnor2_1 _22449_ (.A(_02635_),
    .B(_02642_),
    .Y(_02643_));
 sky130_fd_sc_hd__a21oi_1 _22450_ (.A1(_02630_),
    .A2(_02518_),
    .B1(_02643_),
    .Y(_02644_));
 sky130_fd_sc_hd__and3_1 _22451_ (.A(_02630_),
    .B(_02518_),
    .C(_02643_),
    .X(_02645_));
 sky130_fd_sc_hd__a211o_1 _22452_ (.A1(_02628_),
    .A2(_02629_),
    .B1(_02644_),
    .C1(_02645_),
    .X(_02646_));
 sky130_fd_sc_hd__o211ai_1 _22453_ (.A1(_02644_),
    .A2(_02645_),
    .B1(_02628_),
    .C1(_02629_),
    .Y(_02647_));
 sky130_fd_sc_hd__and2_2 _22454_ (.A(_02646_),
    .B(_02647_),
    .X(_02648_));
 sky130_fd_sc_hd__o21ba_1 _22455_ (.A1(_02521_),
    .A2(_02524_),
    .B1_N(_02522_),
    .X(_02649_));
 sky130_fd_sc_hd__a22oi_2 _22456_ (.A1(_11947_),
    .A2(_12776_),
    .B1(_13960_),
    .B2(_12074_),
    .Y(_02650_));
 sky130_fd_sc_hd__and4_2 _22457_ (.A(_12285_),
    .B(_11830_),
    .C(_13060_),
    .D(_13061_),
    .X(_02651_));
 sky130_fd_sc_hd__o2bb2a_1 _22458_ (.A1_N(_13901_),
    .A2_N(_14499_),
    .B1(_02650_),
    .B2(_02651_),
    .X(_02652_));
 sky130_fd_sc_hd__and4bb_1 _22459_ (.A_N(_02650_),
    .B_N(_02651_),
    .C(_13901_),
    .D(_14324_),
    .X(_02653_));
 sky130_fd_sc_hd__nor2_1 _22460_ (.A(_02652_),
    .B(_02653_),
    .Y(_02654_));
 sky130_fd_sc_hd__xnor2_1 _22461_ (.A(_02649_),
    .B(_02654_),
    .Y(_02655_));
 sky130_fd_sc_hd__o21ai_2 _22462_ (.A1(_02513_),
    .A2(_02515_),
    .B1(_02655_),
    .Y(_02656_));
 sky130_fd_sc_hd__or3_1 _22463_ (.A(_02513_),
    .B(_02515_),
    .C(_02655_),
    .X(_02657_));
 sky130_fd_sc_hd__and2_2 _22464_ (.A(_02656_),
    .B(_02657_),
    .X(_02658_));
 sky130_fd_sc_hd__a22oi_1 _22465_ (.A1(_11825_),
    .A2(_13223_),
    .B1(_14508_),
    .B2(_11482_),
    .Y(_02659_));
 sky130_fd_sc_hd__and4_1 _22466_ (.A(_11834_),
    .B(_11590_),
    .C(_13760_),
    .D(_13545_),
    .X(_02660_));
 sky130_fd_sc_hd__nor2_1 _22467_ (.A(_02659_),
    .B(_02660_),
    .Y(_02661_));
 sky130_fd_sc_hd__nand2_1 _22468_ (.A(_11599_),
    .B(_13054_),
    .Y(_02662_));
 sky130_fd_sc_hd__xnor2_2 _22469_ (.A(_02661_),
    .B(_02662_),
    .Y(_02663_));
 sky130_fd_sc_hd__nand2_1 _22470_ (.A(_11373_),
    .B(_14342_),
    .Y(_02664_));
 sky130_fd_sc_hd__and2b_1 _22471_ (.A_N(_11159_),
    .B(_02237_),
    .X(_02665_));
 sky130_fd_sc_hd__nand2_1 _22472_ (.A(_11171_),
    .B(_14167_),
    .Y(_02666_));
 sky130_fd_sc_hd__xnor2_2 _22473_ (.A(_02665_),
    .B(_02666_),
    .Y(_02667_));
 sky130_fd_sc_hd__xnor2_2 _22474_ (.A(_02664_),
    .B(_02667_),
    .Y(_02668_));
 sky130_fd_sc_hd__and3_1 _22475_ (.A(_11264_),
    .B(_01620_),
    .C(_02527_),
    .X(_02669_));
 sky130_fd_sc_hd__a31o_1 _22476_ (.A1(_11474_),
    .A2(_14343_),
    .A3(_02529_),
    .B1(_02669_),
    .X(_02670_));
 sky130_fd_sc_hd__xor2_2 _22477_ (.A(_02668_),
    .B(_02670_),
    .X(_02671_));
 sky130_fd_sc_hd__xnor2_2 _22478_ (.A(_02663_),
    .B(_02671_),
    .Y(_02672_));
 sky130_fd_sc_hd__nand2_1 _22479_ (.A(_02530_),
    .B(_02532_),
    .Y(_02673_));
 sky130_fd_sc_hd__a21boi_2 _22480_ (.A1(_02525_),
    .A2(_02533_),
    .B1_N(_02673_),
    .Y(_02674_));
 sky130_fd_sc_hd__xnor2_2 _22481_ (.A(_02672_),
    .B(_02674_),
    .Y(_02675_));
 sky130_fd_sc_hd__xnor2_4 _22482_ (.A(_02658_),
    .B(_02675_),
    .Y(_02676_));
 sky130_fd_sc_hd__nand2_1 _22483_ (.A(_02534_),
    .B(_02536_),
    .Y(_02677_));
 sky130_fd_sc_hd__nor2_1 _22484_ (.A(_02534_),
    .B(_02536_),
    .Y(_02678_));
 sky130_fd_sc_hd__a21oi_4 _22485_ (.A1(_02520_),
    .A2(_02677_),
    .B1(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__xnor2_4 _22486_ (.A(_02676_),
    .B(_02679_),
    .Y(_02680_));
 sky130_fd_sc_hd__xnor2_4 _22487_ (.A(_02648_),
    .B(_02680_),
    .Y(_02681_));
 sky130_fd_sc_hd__and2b_1 _22488_ (.A_N(_02541_),
    .B(_02538_),
    .X(_02682_));
 sky130_fd_sc_hd__a21oi_4 _22489_ (.A1(_02510_),
    .A2(_02542_),
    .B1(_02682_),
    .Y(_02683_));
 sky130_fd_sc_hd__xor2_4 _22490_ (.A(_02681_),
    .B(_02683_),
    .X(_02684_));
 sky130_fd_sc_hd__xor2_4 _22491_ (.A(_02627_),
    .B(_02684_),
    .X(_02685_));
 sky130_fd_sc_hd__nor2_1 _22492_ (.A(_02543_),
    .B(_02545_),
    .Y(_02686_));
 sky130_fd_sc_hd__a21oi_2 _22493_ (.A1(_02489_),
    .A2(_02546_),
    .B1(_02686_),
    .Y(_02687_));
 sky130_fd_sc_hd__xnor2_4 _22494_ (.A(_02685_),
    .B(_02687_),
    .Y(_02688_));
 sky130_fd_sc_hd__xnor2_4 _22495_ (.A(_02592_),
    .B(_02688_),
    .Y(_02689_));
 sky130_fd_sc_hd__and2b_1 _22496_ (.A_N(_02549_),
    .B(_02547_),
    .X(_02690_));
 sky130_fd_sc_hd__a21oi_2 _22497_ (.A1(_02455_),
    .A2(_02550_),
    .B1(_02690_),
    .Y(_02691_));
 sky130_fd_sc_hd__xor2_4 _22498_ (.A(_02689_),
    .B(_02691_),
    .X(_02692_));
 sky130_fd_sc_hd__xor2_4 _22499_ (.A(_02572_),
    .B(_02692_),
    .X(_02693_));
 sky130_fd_sc_hd__nor2_1 _22500_ (.A(_02551_),
    .B(_02553_),
    .Y(_02694_));
 sky130_fd_sc_hd__nand2_1 _22501_ (.A(_02551_),
    .B(_02553_),
    .Y(_02695_));
 sky130_fd_sc_hd__o21a_2 _22502_ (.A1(_02432_),
    .A2(_02694_),
    .B1(_02695_),
    .X(_02696_));
 sky130_fd_sc_hd__xnor2_4 _22503_ (.A(_02693_),
    .B(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hd__xnor2_4 _22504_ (.A(_02568_),
    .B(_02697_),
    .Y(_02698_));
 sky130_fd_sc_hd__xor2_4 _22505_ (.A(_02566_),
    .B(_02698_),
    .X(_02699_));
 sky130_fd_sc_hd__or2_1 _22506_ (.A(_02559_),
    .B(_02561_),
    .X(_02700_));
 sky130_fd_sc_hd__a21boi_2 _22507_ (.A1(_02562_),
    .A2(_02564_),
    .B1_N(_02700_),
    .Y(_02701_));
 sky130_fd_sc_hd__xnor2_4 _22508_ (.A(_02699_),
    .B(_02701_),
    .Y(_00089_));
 sky130_fd_sc_hd__a21oi_4 _22509_ (.A1(_02569_),
    .A2(_02570_),
    .B1(_02427_),
    .Y(_02702_));
 sky130_fd_sc_hd__or2b_1 _22510_ (.A(_02574_),
    .B_N(_02590_),
    .X(_02703_));
 sky130_fd_sc_hd__or2b_1 _22511_ (.A(_02573_),
    .B_N(_02591_),
    .X(_02704_));
 sky130_fd_sc_hd__nand2_1 _22512_ (.A(_02703_),
    .B(_02704_),
    .Y(_02705_));
 sky130_fd_sc_hd__xor2_2 _22513_ (.A(_02132_),
    .B(_02705_),
    .X(_02706_));
 sky130_fd_sc_hd__or2b_1 _22514_ (.A(_02588_),
    .B_N(_02585_),
    .X(_02707_));
 sky130_fd_sc_hd__o21a_1 _22515_ (.A1(_02137_),
    .A2(_02589_),
    .B1(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__or3b_1 _22516_ (.A(_02593_),
    .B(_02624_),
    .C_N(_02625_),
    .X(_02709_));
 sky130_fd_sc_hd__and2b_1 _22517_ (.A_N(_02624_),
    .B(_02709_),
    .X(_02710_));
 sky130_fd_sc_hd__or2b_1 _22518_ (.A(_02579_),
    .B_N(_02576_),
    .X(_02711_));
 sky130_fd_sc_hd__a21bo_1 _22519_ (.A1(_02597_),
    .A2(_02605_),
    .B1_N(_02604_),
    .X(_02712_));
 sky130_fd_sc_hd__a31o_1 _22520_ (.A1(_10893_),
    .A2(_13842_),
    .A3(_02595_),
    .B1(_02458_),
    .X(_02713_));
 sky130_fd_sc_hd__xor2_1 _22521_ (.A(_02440_),
    .B(_02713_),
    .X(_02714_));
 sky130_fd_sc_hd__xnor2_1 _22522_ (.A(_02298_),
    .B(_02714_),
    .Y(_02715_));
 sky130_fd_sc_hd__xnor2_1 _22523_ (.A(_02712_),
    .B(_02715_),
    .Y(_02716_));
 sky130_fd_sc_hd__and3_1 _22524_ (.A(_02149_),
    .B(_02151_),
    .C(_02577_),
    .X(_02717_));
 sky130_fd_sc_hd__a21oi_1 _22525_ (.A1(_02445_),
    .A2(_02578_),
    .B1(_02717_),
    .Y(_02718_));
 sky130_fd_sc_hd__xor2_1 _22526_ (.A(_02716_),
    .B(_02718_),
    .X(_02719_));
 sky130_fd_sc_hd__a21oi_1 _22527_ (.A1(_02711_),
    .A2(_02583_),
    .B1(_02719_),
    .Y(_02720_));
 sky130_fd_sc_hd__and3_1 _22528_ (.A(_02711_),
    .B(_02583_),
    .C(_02719_),
    .X(_02721_));
 sky130_fd_sc_hd__nor2_1 _22529_ (.A(_02720_),
    .B(_02721_),
    .Y(_02722_));
 sky130_fd_sc_hd__xnor2_1 _22530_ (.A(_02136_),
    .B(_02722_),
    .Y(_02723_));
 sky130_fd_sc_hd__xnor2_1 _22531_ (.A(_02710_),
    .B(_02723_),
    .Y(_02724_));
 sky130_fd_sc_hd__xnor2_1 _22532_ (.A(_02708_),
    .B(_02724_),
    .Y(_02725_));
 sky130_fd_sc_hd__nor2_1 _22533_ (.A(_02620_),
    .B(_02622_),
    .Y(_02726_));
 sky130_fd_sc_hd__a21o_1 _22534_ (.A1(_02630_),
    .A2(_02518_),
    .B1(_02643_),
    .X(_02727_));
 sky130_fd_sc_hd__nand2_1 _22535_ (.A(_01547_),
    .B(_01846_),
    .Y(_02728_));
 sky130_fd_sc_hd__nand2_1 _22536_ (.A(_11242_),
    .B(_13830_),
    .Y(_02729_));
 sky130_fd_sc_hd__and4_1 _22537_ (.A(_13680_),
    .B(_13678_),
    .C(_13609_),
    .D(_13618_),
    .X(_02730_));
 sky130_fd_sc_hd__a21oi_1 _22538_ (.A1(_02728_),
    .A2(_02729_),
    .B1(_02730_),
    .Y(_02731_));
 sky130_fd_sc_hd__nand2_2 _22539_ (.A(_13897_),
    .B(_14570_),
    .Y(_02732_));
 sky130_fd_sc_hd__xnor2_1 _22540_ (.A(_02731_),
    .B(_02732_),
    .Y(_02733_));
 sky130_fd_sc_hd__nor2_1 _22541_ (.A(_02600_),
    .B(_02602_),
    .Y(_02734_));
 sky130_fd_sc_hd__xnor2_1 _22542_ (.A(_02733_),
    .B(_02734_),
    .Y(_02735_));
 sky130_fd_sc_hd__nand2_1 _22543_ (.A(_02598_),
    .B(_02735_),
    .Y(_02736_));
 sky130_fd_sc_hd__or2_1 _22544_ (.A(_02597_),
    .B(_02735_),
    .X(_02737_));
 sky130_fd_sc_hd__nand2_1 _22545_ (.A(_02736_),
    .B(_02737_),
    .Y(_02738_));
 sky130_fd_sc_hd__or2b_1 _22546_ (.A(_02612_),
    .B_N(_02617_),
    .X(_02739_));
 sky130_fd_sc_hd__nand2_1 _22547_ (.A(_02611_),
    .B(_02618_),
    .Y(_02740_));
 sky130_fd_sc_hd__a31o_1 _22548_ (.A1(_14099_),
    .A2(_01718_),
    .A3(_02615_),
    .B1(_02614_),
    .X(_02741_));
 sky130_fd_sc_hd__o21ba_1 _22549_ (.A1(_02631_),
    .A2(_02634_),
    .B1_N(_02632_),
    .X(_02742_));
 sky130_fd_sc_hd__a22oi_1 _22550_ (.A1(_11927_),
    .A2(_14417_),
    .B1(_13839_),
    .B2(_14105_),
    .Y(_02743_));
 sky130_fd_sc_hd__and4_1 _22551_ (.A(_14103_),
    .B(_13691_),
    .C(_13445_),
    .D(_13281_),
    .X(_02744_));
 sky130_fd_sc_hd__nor2_1 _22552_ (.A(_02743_),
    .B(_02744_),
    .Y(_02745_));
 sky130_fd_sc_hd__nand2_1 _22553_ (.A(_11775_),
    .B(_13824_),
    .Y(_02746_));
 sky130_fd_sc_hd__xnor2_2 _22554_ (.A(_02745_),
    .B(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__xnor2_1 _22555_ (.A(_02742_),
    .B(_02747_),
    .Y(_02748_));
 sky130_fd_sc_hd__xnor2_1 _22556_ (.A(_02741_),
    .B(_02748_),
    .Y(_02749_));
 sky130_fd_sc_hd__a21oi_1 _22557_ (.A1(_02739_),
    .A2(_02740_),
    .B1(_02749_),
    .Y(_02750_));
 sky130_fd_sc_hd__and3_1 _22558_ (.A(_02739_),
    .B(_02740_),
    .C(_02749_),
    .X(_02751_));
 sky130_fd_sc_hd__nor3_1 _22559_ (.A(_02738_),
    .B(_02750_),
    .C(_02751_),
    .Y(_02752_));
 sky130_fd_sc_hd__o21a_1 _22560_ (.A1(_02750_),
    .A2(_02751_),
    .B1(_02738_),
    .X(_02753_));
 sky130_fd_sc_hd__a211oi_1 _22561_ (.A1(_02727_),
    .A2(_02646_),
    .B1(_02752_),
    .C1(_02753_),
    .Y(_02754_));
 sky130_fd_sc_hd__o211ai_1 _22562_ (.A1(_02752_),
    .A2(_02753_),
    .B1(_02727_),
    .C1(_02646_),
    .Y(_02755_));
 sky130_fd_sc_hd__and2b_1 _22563_ (.A_N(_02754_),
    .B(_02755_),
    .X(_02756_));
 sky130_fd_sc_hd__xnor2_1 _22564_ (.A(_02726_),
    .B(_02756_),
    .Y(_02757_));
 sky130_fd_sc_hd__or2b_1 _22565_ (.A(_02641_),
    .B_N(_02640_),
    .X(_02758_));
 sky130_fd_sc_hd__nand2_1 _22566_ (.A(_02635_),
    .B(_02642_),
    .Y(_02759_));
 sky130_fd_sc_hd__or3_1 _22567_ (.A(_02649_),
    .B(_02652_),
    .C(_02653_),
    .X(_02760_));
 sky130_fd_sc_hd__a22oi_2 _22568_ (.A1(_13716_),
    .A2(_14076_),
    .B1(_13637_),
    .B2(_11891_),
    .Y(_02761_));
 sky130_fd_sc_hd__and4_1 _22569_ (.A(_14123_),
    .B(_12023_),
    .C(_13859_),
    .D(_13125_),
    .X(_02762_));
 sky130_fd_sc_hd__nor2_1 _22570_ (.A(_02761_),
    .B(_02762_),
    .Y(_02763_));
 sky130_fd_sc_hd__nand2_1 _22571_ (.A(_12591_),
    .B(_13868_),
    .Y(_02764_));
 sky130_fd_sc_hd__xnor2_1 _22572_ (.A(_02763_),
    .B(_02764_),
    .Y(_02765_));
 sky130_fd_sc_hd__a22oi_2 _22573_ (.A1(_14131_),
    .A2(_12983_),
    .B1(_13944_),
    .B2(_12271_),
    .Y(_02766_));
 sky130_fd_sc_hd__and4_1 _22574_ (.A(_12273_),
    .B(_12328_),
    .C(_12983_),
    .D(_13376_),
    .X(_02767_));
 sky130_fd_sc_hd__nor2_1 _22575_ (.A(_02766_),
    .B(_02767_),
    .Y(_02768_));
 sky130_fd_sc_hd__nand2_1 _22576_ (.A(_12226_),
    .B(_14080_),
    .Y(_02769_));
 sky130_fd_sc_hd__xnor2_1 _22577_ (.A(_02768_),
    .B(_02769_),
    .Y(_02770_));
 sky130_fd_sc_hd__o21ba_1 _22578_ (.A1(_02636_),
    .A2(_02639_),
    .B1_N(_02637_),
    .X(_02771_));
 sky130_fd_sc_hd__xnor2_1 _22579_ (.A(_02770_),
    .B(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__xnor2_1 _22580_ (.A(_02765_),
    .B(_02772_),
    .Y(_02773_));
 sky130_fd_sc_hd__a21oi_1 _22581_ (.A1(_02760_),
    .A2(_02656_),
    .B1(_02773_),
    .Y(_02774_));
 sky130_fd_sc_hd__and3_1 _22582_ (.A(_02760_),
    .B(_02656_),
    .C(_02773_),
    .X(_02775_));
 sky130_fd_sc_hd__a211o_1 _22583_ (.A1(_02758_),
    .A2(_02759_),
    .B1(_02774_),
    .C1(_02775_),
    .X(_02776_));
 sky130_fd_sc_hd__o211ai_1 _22584_ (.A1(_02774_),
    .A2(_02775_),
    .B1(_02758_),
    .C1(_02759_),
    .Y(_02777_));
 sky130_fd_sc_hd__and2_1 _22585_ (.A(_02776_),
    .B(_02777_),
    .X(_02778_));
 sky130_fd_sc_hd__o21ba_1 _22586_ (.A1(_02659_),
    .A2(_02662_),
    .B1_N(_02660_),
    .X(_02779_));
 sky130_fd_sc_hd__a22oi_1 _22587_ (.A1(_13305_),
    .A2(_13555_),
    .B1(_01601_),
    .B2(_11949_),
    .Y(_02780_));
 sky130_fd_sc_hd__and4_2 _22588_ (.A(_11946_),
    .B(_11958_),
    .C(_12770_),
    .D(_12910_),
    .X(_02781_));
 sky130_fd_sc_hd__o2bb2a_1 _22589_ (.A1_N(_13666_),
    .A2_N(_14324_),
    .B1(_02780_),
    .B2(_02781_),
    .X(_02782_));
 sky130_fd_sc_hd__and4bb_2 _22590_ (.A_N(_02780_),
    .B_N(_02781_),
    .C(_12145_),
    .D(_12584_),
    .X(_02783_));
 sky130_fd_sc_hd__nor2_1 _22591_ (.A(_02782_),
    .B(_02783_),
    .Y(_02784_));
 sky130_fd_sc_hd__xnor2_1 _22592_ (.A(_02779_),
    .B(_02784_),
    .Y(_02785_));
 sky130_fd_sc_hd__o21ai_2 _22593_ (.A1(_02651_),
    .A2(_02653_),
    .B1(_02785_),
    .Y(_02786_));
 sky130_fd_sc_hd__or3_1 _22594_ (.A(_02651_),
    .B(_02653_),
    .C(_02785_),
    .X(_02787_));
 sky130_fd_sc_hd__and2_1 _22595_ (.A(_02786_),
    .B(_02787_),
    .X(_02788_));
 sky130_fd_sc_hd__a22oi_1 _22596_ (.A1(_13695_),
    .A2(_13228_),
    .B1(_13762_),
    .B2(_11591_),
    .Y(_02789_));
 sky130_fd_sc_hd__and4_1 _22597_ (.A(_11490_),
    .B(_11699_),
    .C(_13223_),
    .D(_13971_),
    .X(_02790_));
 sky130_fd_sc_hd__nor2_1 _22598_ (.A(_02789_),
    .B(_02790_),
    .Y(_02791_));
 sky130_fd_sc_hd__nand2_1 _22599_ (.A(_11820_),
    .B(_14154_),
    .Y(_02792_));
 sky130_fd_sc_hd__xnor2_2 _22600_ (.A(_02791_),
    .B(_02792_),
    .Y(_02793_));
 sky130_fd_sc_hd__nand2_1 _22601_ (.A(_11482_),
    .B(\genblk1.pcpi_mul.rs2[30] ),
    .Y(_02794_));
 sky130_fd_sc_hd__and2b_1 _22602_ (.A_N(_12098_),
    .B(\genblk1.pcpi_mul.rs2[32] ),
    .X(_02795_));
 sky130_fd_sc_hd__nand2_1 _22603_ (.A(_11712_),
    .B(\genblk1.pcpi_mul.rs2[31] ),
    .Y(_02796_));
 sky130_fd_sc_hd__xnor2_2 _22604_ (.A(_02795_),
    .B(_02796_),
    .Y(_02797_));
 sky130_fd_sc_hd__xnor2_2 _22605_ (.A(_02794_),
    .B(_02797_),
    .Y(_02798_));
 sky130_fd_sc_hd__and3_1 _22606_ (.A(_11261_),
    .B(_13753_),
    .C(_02665_),
    .X(_02799_));
 sky130_fd_sc_hd__a31o_1 _22607_ (.A1(_11278_),
    .A2(_14160_),
    .A3(_02667_),
    .B1(_02799_),
    .X(_02800_));
 sky130_fd_sc_hd__xor2_2 _22608_ (.A(_02798_),
    .B(_02800_),
    .X(_02801_));
 sky130_fd_sc_hd__xnor2_2 _22609_ (.A(_02793_),
    .B(_02801_),
    .Y(_02802_));
 sky130_fd_sc_hd__nand2_1 _22610_ (.A(_02668_),
    .B(_02670_),
    .Y(_02803_));
 sky130_fd_sc_hd__a21boi_2 _22611_ (.A1(_02663_),
    .A2(_02671_),
    .B1_N(_02803_),
    .Y(_02804_));
 sky130_fd_sc_hd__xnor2_1 _22612_ (.A(_02802_),
    .B(_02804_),
    .Y(_02805_));
 sky130_fd_sc_hd__xnor2_2 _22613_ (.A(_02788_),
    .B(_02805_),
    .Y(_02806_));
 sky130_fd_sc_hd__nand2_1 _22614_ (.A(_02672_),
    .B(_02674_),
    .Y(_02807_));
 sky130_fd_sc_hd__nor2_1 _22615_ (.A(_02672_),
    .B(_02674_),
    .Y(_02808_));
 sky130_fd_sc_hd__a21oi_2 _22616_ (.A1(_02658_),
    .A2(_02807_),
    .B1(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hd__xnor2_2 _22617_ (.A(_02806_),
    .B(_02809_),
    .Y(_02810_));
 sky130_fd_sc_hd__xnor2_2 _22618_ (.A(_02778_),
    .B(_02810_),
    .Y(_02811_));
 sky130_fd_sc_hd__and2b_1 _22619_ (.A_N(_02679_),
    .B(_02676_),
    .X(_02812_));
 sky130_fd_sc_hd__a21oi_2 _22620_ (.A1(_02648_),
    .A2(_02680_),
    .B1(_02812_),
    .Y(_02813_));
 sky130_fd_sc_hd__xor2_1 _22621_ (.A(_02811_),
    .B(_02813_),
    .X(_02814_));
 sky130_fd_sc_hd__xor2_1 _22622_ (.A(_02757_),
    .B(_02814_),
    .X(_02815_));
 sky130_fd_sc_hd__nor2_1 _22623_ (.A(_02681_),
    .B(_02683_),
    .Y(_02816_));
 sky130_fd_sc_hd__a21oi_1 _22624_ (.A1(_02627_),
    .A2(_02684_),
    .B1(_02816_),
    .Y(_02817_));
 sky130_fd_sc_hd__xnor2_1 _22625_ (.A(_02815_),
    .B(_02817_),
    .Y(_02818_));
 sky130_fd_sc_hd__xor2_1 _22626_ (.A(_02725_),
    .B(_02818_),
    .X(_02819_));
 sky130_fd_sc_hd__and2b_1 _22627_ (.A_N(_02687_),
    .B(_02685_),
    .X(_02820_));
 sky130_fd_sc_hd__a21o_1 _22628_ (.A1(_02592_),
    .A2(_02688_),
    .B1(_02820_),
    .X(_02821_));
 sky130_fd_sc_hd__xor2_1 _22629_ (.A(_02819_),
    .B(_02821_),
    .X(_02822_));
 sky130_fd_sc_hd__xnor2_2 _22630_ (.A(_02706_),
    .B(_02822_),
    .Y(_02823_));
 sky130_fd_sc_hd__nor2_1 _22631_ (.A(_02689_),
    .B(_02691_),
    .Y(_02824_));
 sky130_fd_sc_hd__a21oi_2 _22632_ (.A1(_02572_),
    .A2(_02692_),
    .B1(_02824_),
    .Y(_02825_));
 sky130_fd_sc_hd__xnor2_2 _22633_ (.A(_02823_),
    .B(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__xnor2_4 _22634_ (.A(_02702_),
    .B(_02826_),
    .Y(_02827_));
 sky130_fd_sc_hd__or2b_1 _22635_ (.A(_02696_),
    .B_N(_02693_),
    .X(_02828_));
 sky130_fd_sc_hd__a21boi_4 _22636_ (.A1(_02568_),
    .A2(_02697_),
    .B1_N(_02828_),
    .Y(_02829_));
 sky130_fd_sc_hd__xnor2_4 _22637_ (.A(_02827_),
    .B(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__nand2_1 _22638_ (.A(_02562_),
    .B(_02699_),
    .Y(_02831_));
 sky130_vsdinv _22639_ (.A(_02831_),
    .Y(_02832_));
 sky130_fd_sc_hd__o21a_1 _22640_ (.A1(_02566_),
    .A2(_02698_),
    .B1(_02700_),
    .X(_02833_));
 sky130_fd_sc_hd__a21o_1 _22641_ (.A1(_02566_),
    .A2(_02698_),
    .B1(_02833_),
    .X(_02834_));
 sky130_fd_sc_hd__a21boi_4 _22642_ (.A1(_02564_),
    .A2(_02832_),
    .B1_N(_02834_),
    .Y(_02835_));
 sky130_fd_sc_hd__xor2_4 _22643_ (.A(_02830_),
    .B(_02835_),
    .X(_00090_));
 sky130_fd_sc_hd__or2b_1 _22644_ (.A(_02825_),
    .B_N(_02823_),
    .X(_02836_));
 sky130_fd_sc_hd__nand2_1 _22645_ (.A(_02702_),
    .B(_02826_),
    .Y(_02837_));
 sky130_fd_sc_hd__a21oi_1 _22646_ (.A1(_02703_),
    .A2(_02704_),
    .B1(_02427_),
    .Y(_02838_));
 sky130_fd_sc_hd__or2b_1 _22647_ (.A(_02710_),
    .B_N(_02723_),
    .X(_02839_));
 sky130_fd_sc_hd__or2b_1 _22648_ (.A(_02708_),
    .B_N(_02724_),
    .X(_02840_));
 sky130_fd_sc_hd__nand2_1 _22649_ (.A(_02839_),
    .B(_02840_),
    .Y(_02841_));
 sky130_fd_sc_hd__xor2_1 _22650_ (.A(_02287_),
    .B(_02841_),
    .X(_02842_));
 sky130_fd_sc_hd__and2b_1 _22651_ (.A_N(_02137_),
    .B(_02722_),
    .X(_02843_));
 sky130_fd_sc_hd__nor2_1 _22652_ (.A(_02720_),
    .B(_02843_),
    .Y(_02844_));
 sky130_fd_sc_hd__or3b_1 _22653_ (.A(_02726_),
    .B(_02754_),
    .C_N(_02755_),
    .X(_02845_));
 sky130_fd_sc_hd__and2b_1 _22654_ (.A_N(_02754_),
    .B(_02845_),
    .X(_02846_));
 sky130_fd_sc_hd__or2b_1 _22655_ (.A(_02734_),
    .B_N(_02733_),
    .X(_02847_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _22656_ (.A(_02715_),
    .X(_02848_));
 sky130_fd_sc_hd__a21o_1 _22657_ (.A1(_02847_),
    .A2(_02736_),
    .B1(_02848_),
    .X(_02849_));
 sky130_fd_sc_hd__nand3_1 _22658_ (.A(_02848_),
    .B(_02847_),
    .C(_02736_),
    .Y(_02850_));
 sky130_fd_sc_hd__nand2_1 _22659_ (.A(_02849_),
    .B(_02850_),
    .Y(_02851_));
 sky130_fd_sc_hd__or2_1 _22660_ (.A(_02440_),
    .B(_02713_),
    .X(_02852_));
 sky130_fd_sc_hd__and3_1 _22661_ (.A(_02149_),
    .B(_02151_),
    .C(_02713_),
    .X(_02853_));
 sky130_fd_sc_hd__a21oi_4 _22662_ (.A1(_02445_),
    .A2(_02852_),
    .B1(_02853_),
    .Y(_02854_));
 sky130_fd_sc_hd__xnor2_1 _22663_ (.A(_02851_),
    .B(_02854_),
    .Y(_02855_));
 sky130_fd_sc_hd__or2b_1 _22664_ (.A(_02848_),
    .B_N(_02712_),
    .X(_02856_));
 sky130_fd_sc_hd__or2b_1 _22665_ (.A(_02718_),
    .B_N(_02716_),
    .X(_02857_));
 sky130_fd_sc_hd__nand2_1 _22666_ (.A(_02856_),
    .B(_02857_),
    .Y(_02858_));
 sky130_fd_sc_hd__xor2_1 _22667_ (.A(_02855_),
    .B(_02858_),
    .X(_02859_));
 sky130_fd_sc_hd__xor2_1 _22668_ (.A(_01995_),
    .B(_02859_),
    .X(_02860_));
 sky130_fd_sc_hd__xnor2_1 _22669_ (.A(_02846_),
    .B(_02860_),
    .Y(_02861_));
 sky130_fd_sc_hd__xnor2_1 _22670_ (.A(_02844_),
    .B(_02861_),
    .Y(_02862_));
 sky130_fd_sc_hd__nor2_1 _22671_ (.A(_02750_),
    .B(_02752_),
    .Y(_02863_));
 sky130_fd_sc_hd__a21o_1 _22672_ (.A1(_02760_),
    .A2(_02656_),
    .B1(_02773_),
    .X(_02864_));
 sky130_fd_sc_hd__a31oi_2 _22673_ (.A1(_11137_),
    .A2(_14562_),
    .A3(_02731_),
    .B1(_02730_),
    .Y(_02865_));
 sky130_fd_sc_hd__nand2_1 _22674_ (.A(_01547_),
    .B(_14026_),
    .Y(_02866_));
 sky130_fd_sc_hd__a22o_1 _22675_ (.A1(_13900_),
    .A2(_13618_),
    .B1(_13842_),
    .B2(_13899_),
    .X(_02867_));
 sky130_fd_sc_hd__o21a_1 _22676_ (.A1(_02729_),
    .A2(_02866_),
    .B1(_02867_),
    .X(_02868_));
 sky130_fd_sc_hd__xnor2_1 _22677_ (.A(_02732_),
    .B(_02868_),
    .Y(_02869_));
 sky130_fd_sc_hd__xnor2_1 _22678_ (.A(_02865_),
    .B(_02869_),
    .Y(_02870_));
 sky130_fd_sc_hd__nand2_1 _22679_ (.A(_02597_),
    .B(_02870_),
    .Y(_02871_));
 sky130_fd_sc_hd__or2_1 _22680_ (.A(_02597_),
    .B(_02870_),
    .X(_02872_));
 sky130_fd_sc_hd__nand2_1 _22681_ (.A(_02871_),
    .B(_02872_),
    .Y(_02873_));
 sky130_fd_sc_hd__or2b_1 _22682_ (.A(_02742_),
    .B_N(_02747_),
    .X(_02874_));
 sky130_fd_sc_hd__nand2_1 _22683_ (.A(_02741_),
    .B(_02748_),
    .Y(_02875_));
 sky130_fd_sc_hd__a31o_1 _22684_ (.A1(_14099_),
    .A2(_13815_),
    .A3(_02745_),
    .B1(_02744_),
    .X(_02876_));
 sky130_fd_sc_hd__o21ba_1 _22685_ (.A1(_02761_),
    .A2(_02764_),
    .B1_N(_02762_),
    .X(_02877_));
 sky130_fd_sc_hd__a22oi_1 _22686_ (.A1(_11665_),
    .A2(_14418_),
    .B1(_13813_),
    .B2(_11556_),
    .Y(_02878_));
 sky130_fd_sc_hd__and4_1 _22687_ (.A(_11663_),
    .B(_11925_),
    .C(_13128_),
    .D(_13292_),
    .X(_02879_));
 sky130_fd_sc_hd__nor2_1 _22688_ (.A(_02878_),
    .B(_02879_),
    .Y(_02880_));
 sky130_fd_sc_hd__nand2_1 _22689_ (.A(_11560_),
    .B(_14225_),
    .Y(_02881_));
 sky130_fd_sc_hd__xnor2_1 _22690_ (.A(_02880_),
    .B(_02881_),
    .Y(_02882_));
 sky130_fd_sc_hd__xnor2_1 _22691_ (.A(_02877_),
    .B(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__xnor2_1 _22692_ (.A(_02876_),
    .B(_02883_),
    .Y(_02884_));
 sky130_fd_sc_hd__a21oi_1 _22693_ (.A1(_02874_),
    .A2(_02875_),
    .B1(_02884_),
    .Y(_02885_));
 sky130_fd_sc_hd__and3_1 _22694_ (.A(_02874_),
    .B(_02875_),
    .C(_02884_),
    .X(_02886_));
 sky130_fd_sc_hd__nor3_1 _22695_ (.A(_02873_),
    .B(_02885_),
    .C(_02886_),
    .Y(_02887_));
 sky130_fd_sc_hd__o21a_1 _22696_ (.A1(_02885_),
    .A2(_02886_),
    .B1(_02873_),
    .X(_02888_));
 sky130_fd_sc_hd__a211oi_1 _22697_ (.A1(_02864_),
    .A2(_02776_),
    .B1(_02887_),
    .C1(_02888_),
    .Y(_02889_));
 sky130_fd_sc_hd__o211ai_1 _22698_ (.A1(_02887_),
    .A2(_02888_),
    .B1(_02864_),
    .C1(_02776_),
    .Y(_02890_));
 sky130_fd_sc_hd__and2b_1 _22699_ (.A_N(_02889_),
    .B(_02890_),
    .X(_02891_));
 sky130_fd_sc_hd__xnor2_1 _22700_ (.A(_02863_),
    .B(_02891_),
    .Y(_02892_));
 sky130_fd_sc_hd__or2b_1 _22701_ (.A(_02771_),
    .B_N(_02770_),
    .X(_02893_));
 sky130_fd_sc_hd__nand2_1 _22702_ (.A(_02765_),
    .B(_02772_),
    .Y(_02894_));
 sky130_fd_sc_hd__or3_2 _22703_ (.A(_02779_),
    .B(_02782_),
    .C(_02783_),
    .X(_02895_));
 sky130_fd_sc_hd__a22oi_1 _22704_ (.A1(_12023_),
    .A2(_13125_),
    .B1(_14056_),
    .B2(_14123_),
    .Y(_02896_));
 sky130_fd_sc_hd__and4_1 _22705_ (.A(_11890_),
    .B(_13715_),
    .C(_13636_),
    .D(_13867_),
    .X(_02897_));
 sky130_fd_sc_hd__nor2_1 _22706_ (.A(_02896_),
    .B(_02897_),
    .Y(_02898_));
 sky130_fd_sc_hd__nand2_1 _22707_ (.A(_12591_),
    .B(_13838_),
    .Y(_02899_));
 sky130_fd_sc_hd__xnor2_2 _22708_ (.A(_02898_),
    .B(_02899_),
    .Y(_02900_));
 sky130_fd_sc_hd__a22oi_1 _22709_ (.A1(_14268_),
    .A2(_14129_),
    .B1(_12830_),
    .B2(_12329_),
    .Y(_02901_));
 sky130_fd_sc_hd__and4_1 _22710_ (.A(_01912_),
    .B(_12282_),
    .C(_13944_),
    .D(_12416_),
    .X(_02902_));
 sky130_fd_sc_hd__nor2_1 _22711_ (.A(_02901_),
    .B(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__nand2_1 _22712_ (.A(_12227_),
    .B(_13860_),
    .Y(_02904_));
 sky130_fd_sc_hd__xnor2_2 _22713_ (.A(_02903_),
    .B(_02904_),
    .Y(_02905_));
 sky130_fd_sc_hd__o21ba_1 _22714_ (.A1(_02766_),
    .A2(_02769_),
    .B1_N(_02767_),
    .X(_02906_));
 sky130_fd_sc_hd__xnor2_2 _22715_ (.A(_02905_),
    .B(_02906_),
    .Y(_02907_));
 sky130_fd_sc_hd__xnor2_2 _22716_ (.A(_02900_),
    .B(_02907_),
    .Y(_02908_));
 sky130_fd_sc_hd__a21oi_4 _22717_ (.A1(_02895_),
    .A2(_02786_),
    .B1(_02908_),
    .Y(_02909_));
 sky130_fd_sc_hd__and3_1 _22718_ (.A(_02895_),
    .B(_02786_),
    .C(_02908_),
    .X(_02910_));
 sky130_fd_sc_hd__a211oi_4 _22719_ (.A1(_02893_),
    .A2(_02894_),
    .B1(_02909_),
    .C1(_02910_),
    .Y(_02911_));
 sky130_fd_sc_hd__o211a_1 _22720_ (.A1(_02909_),
    .A2(_02910_),
    .B1(_02893_),
    .C1(_02894_),
    .X(_02912_));
 sky130_fd_sc_hd__nor2_2 _22721_ (.A(_02911_),
    .B(_02912_),
    .Y(_02913_));
 sky130_fd_sc_hd__o21ba_1 _22722_ (.A1(_02789_),
    .A2(_02792_),
    .B1_N(_02790_),
    .X(_02914_));
 sky130_fd_sc_hd__a22oi_1 _22723_ (.A1(_12079_),
    .A2(_12771_),
    .B1(_13960_),
    .B2(_12070_),
    .Y(_02915_));
 sky130_fd_sc_hd__and4_2 _22724_ (.A(_12067_),
    .B(_12144_),
    .C(_13558_),
    .D(_13740_),
    .X(_02916_));
 sky130_fd_sc_hd__o2bb2a_1 _22725_ (.A1_N(_13484_),
    .A2_N(_14499_),
    .B1(_02915_),
    .B2(_02916_),
    .X(_02917_));
 sky130_fd_sc_hd__and4bb_2 _22726_ (.A_N(_02915_),
    .B_N(_02916_),
    .C(_14272_),
    .D(_14324_),
    .X(_02918_));
 sky130_fd_sc_hd__nor2_1 _22727_ (.A(_02917_),
    .B(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__xnor2_2 _22728_ (.A(_02914_),
    .B(_02919_),
    .Y(_02920_));
 sky130_fd_sc_hd__o21ai_4 _22729_ (.A1(_02781_),
    .A2(_02783_),
    .B1(_02920_),
    .Y(_02921_));
 sky130_fd_sc_hd__or3_1 _22730_ (.A(_02781_),
    .B(_02783_),
    .C(_02920_),
    .X(_02922_));
 sky130_fd_sc_hd__and2_2 _22731_ (.A(_02921_),
    .B(_02922_),
    .X(_02923_));
 sky130_fd_sc_hd__a22oi_2 _22732_ (.A1(_13918_),
    .A2(_13764_),
    .B1(_14508_),
    .B2(_11599_),
    .Y(_02924_));
 sky130_fd_sc_hd__and4_1 _22733_ (.A(_13689_),
    .B(_12074_),
    .C(_13760_),
    .D(_13545_),
    .X(_02925_));
 sky130_fd_sc_hd__nor2_1 _22734_ (.A(_02924_),
    .B(_02925_),
    .Y(_02926_));
 sky130_fd_sc_hd__nand2_1 _22735_ (.A(_11950_),
    .B(_14154_),
    .Y(_02927_));
 sky130_fd_sc_hd__xnor2_2 _22736_ (.A(_02926_),
    .B(_02927_),
    .Y(_02928_));
 sky130_fd_sc_hd__nand2_1 _22737_ (.A(_11591_),
    .B(_13541_),
    .Y(_02929_));
 sky130_fd_sc_hd__and2b_1 _22738_ (.A_N(_11276_),
    .B(_02237_),
    .X(_02930_));
 sky130_fd_sc_hd__nand2_1 _22739_ (.A(_11380_),
    .B(_14167_),
    .Y(_02931_));
 sky130_fd_sc_hd__xnor2_2 _22740_ (.A(_02930_),
    .B(_02931_),
    .Y(_02932_));
 sky130_fd_sc_hd__xnor2_2 _22741_ (.A(_02929_),
    .B(_02932_),
    .Y(_02933_));
 sky130_fd_sc_hd__and3_1 _22742_ (.A(_12343_),
    .B(_01620_),
    .C(_02795_),
    .X(_02934_));
 sky130_fd_sc_hd__a31o_1 _22743_ (.A1(_11382_),
    .A2(_14343_),
    .A3(_02797_),
    .B1(_02934_),
    .X(_02935_));
 sky130_fd_sc_hd__xor2_2 _22744_ (.A(_02933_),
    .B(_02935_),
    .X(_02936_));
 sky130_fd_sc_hd__xnor2_2 _22745_ (.A(_02928_),
    .B(_02936_),
    .Y(_02937_));
 sky130_fd_sc_hd__nand2_1 _22746_ (.A(_02798_),
    .B(_02800_),
    .Y(_02938_));
 sky130_fd_sc_hd__a21boi_2 _22747_ (.A1(_02793_),
    .A2(_02801_),
    .B1_N(_02938_),
    .Y(_02939_));
 sky130_fd_sc_hd__xnor2_1 _22748_ (.A(_02937_),
    .B(_02939_),
    .Y(_02940_));
 sky130_fd_sc_hd__xnor2_2 _22749_ (.A(_02923_),
    .B(_02940_),
    .Y(_02941_));
 sky130_fd_sc_hd__nand2_1 _22750_ (.A(_02802_),
    .B(_02804_),
    .Y(_02942_));
 sky130_fd_sc_hd__nor2_1 _22751_ (.A(_02802_),
    .B(_02804_),
    .Y(_02943_));
 sky130_fd_sc_hd__a21oi_2 _22752_ (.A1(_02788_),
    .A2(_02942_),
    .B1(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__xnor2_2 _22753_ (.A(_02941_),
    .B(_02944_),
    .Y(_02945_));
 sky130_fd_sc_hd__xnor2_2 _22754_ (.A(_02913_),
    .B(_02945_),
    .Y(_02946_));
 sky130_fd_sc_hd__and2b_1 _22755_ (.A_N(_02809_),
    .B(_02806_),
    .X(_02947_));
 sky130_fd_sc_hd__a21oi_2 _22756_ (.A1(_02778_),
    .A2(_02810_),
    .B1(_02947_),
    .Y(_02948_));
 sky130_fd_sc_hd__xor2_1 _22757_ (.A(_02946_),
    .B(_02948_),
    .X(_02949_));
 sky130_fd_sc_hd__xor2_1 _22758_ (.A(_02892_),
    .B(_02949_),
    .X(_02950_));
 sky130_fd_sc_hd__nor2_1 _22759_ (.A(_02811_),
    .B(_02813_),
    .Y(_02951_));
 sky130_fd_sc_hd__a21oi_1 _22760_ (.A1(_02757_),
    .A2(_02814_),
    .B1(_02951_),
    .Y(_02952_));
 sky130_fd_sc_hd__xnor2_1 _22761_ (.A(_02950_),
    .B(_02952_),
    .Y(_02953_));
 sky130_fd_sc_hd__xor2_1 _22762_ (.A(_02862_),
    .B(_02953_),
    .X(_02954_));
 sky130_fd_sc_hd__and2b_1 _22763_ (.A_N(_02817_),
    .B(_02815_),
    .X(_02955_));
 sky130_fd_sc_hd__a21o_1 _22764_ (.A1(_02725_),
    .A2(_02818_),
    .B1(_02955_),
    .X(_02956_));
 sky130_fd_sc_hd__xor2_1 _22765_ (.A(_02954_),
    .B(_02956_),
    .X(_02957_));
 sky130_fd_sc_hd__xnor2_1 _22766_ (.A(_02842_),
    .B(_02957_),
    .Y(_02958_));
 sky130_fd_sc_hd__nor2_1 _22767_ (.A(_02819_),
    .B(_02821_),
    .Y(_02959_));
 sky130_fd_sc_hd__nand2_1 _22768_ (.A(_02819_),
    .B(_02821_),
    .Y(_02960_));
 sky130_fd_sc_hd__o21a_1 _22769_ (.A1(_02706_),
    .A2(_02959_),
    .B1(_02960_),
    .X(_02961_));
 sky130_fd_sc_hd__xnor2_1 _22770_ (.A(_02958_),
    .B(_02961_),
    .Y(_02962_));
 sky130_fd_sc_hd__xnor2_1 _22771_ (.A(_02838_),
    .B(_02962_),
    .Y(_02963_));
 sky130_fd_sc_hd__a21o_1 _22772_ (.A1(_02836_),
    .A2(_02837_),
    .B1(_02963_),
    .X(_02964_));
 sky130_vsdinv _22773_ (.A(_02964_),
    .Y(_02965_));
 sky130_fd_sc_hd__and3_1 _22774_ (.A(_02836_),
    .B(_02837_),
    .C(_02963_),
    .X(_02966_));
 sky130_fd_sc_hd__nor2_2 _22775_ (.A(_02965_),
    .B(_02966_),
    .Y(_02967_));
 sky130_fd_sc_hd__or2_1 _22776_ (.A(_02827_),
    .B(_02829_),
    .X(_02968_));
 sky130_fd_sc_hd__o21ai_2 _22777_ (.A1(_02830_),
    .A2(_02835_),
    .B1(_02968_),
    .Y(_02969_));
 sky130_fd_sc_hd__xor2_4 _22778_ (.A(_02967_),
    .B(_02969_),
    .X(_00091_));
 sky130_fd_sc_hd__a21oi_4 _22779_ (.A1(_02839_),
    .A2(_02840_),
    .B1(_02427_),
    .Y(_02970_));
 sky130_fd_sc_hd__or2b_1 _22780_ (.A(_02846_),
    .B_N(_02860_),
    .X(_02971_));
 sky130_fd_sc_hd__or2b_1 _22781_ (.A(_02844_),
    .B_N(_02861_),
    .X(_02972_));
 sky130_fd_sc_hd__nand2_1 _22782_ (.A(_02971_),
    .B(_02972_),
    .Y(_02973_));
 sky130_fd_sc_hd__xor2_2 _22783_ (.A(_02287_),
    .B(_02973_),
    .X(_02974_));
 sky130_fd_sc_hd__or2b_1 _22784_ (.A(_02855_),
    .B_N(_02858_),
    .X(_02975_));
 sky130_fd_sc_hd__o21ai_1 _22785_ (.A1(_02433_),
    .A2(_02859_),
    .B1(_02975_),
    .Y(_02976_));
 sky130_fd_sc_hd__or3b_1 _22786_ (.A(_02863_),
    .B(_02889_),
    .C_N(_02890_),
    .X(_02977_));
 sky130_fd_sc_hd__and2b_1 _22787_ (.A_N(_02889_),
    .B(_02977_),
    .X(_02978_));
 sky130_fd_sc_hd__or2b_1 _22788_ (.A(_02865_),
    .B_N(_02869_),
    .X(_02979_));
 sky130_fd_sc_hd__a21o_1 _22789_ (.A1(_02979_),
    .A2(_02871_),
    .B1(_02848_),
    .X(_02980_));
 sky130_fd_sc_hd__nand3_1 _22790_ (.A(_02848_),
    .B(_02979_),
    .C(_02871_),
    .Y(_02981_));
 sky130_fd_sc_hd__nand2_1 _22791_ (.A(_02980_),
    .B(_02981_),
    .Y(_02982_));
 sky130_fd_sc_hd__xor2_1 _22792_ (.A(_02854_),
    .B(_02982_),
    .X(_02983_));
 sky130_fd_sc_hd__o21a_1 _22793_ (.A1(_02851_),
    .A2(_02854_),
    .B1(_02849_),
    .X(_02984_));
 sky130_fd_sc_hd__xor2_1 _22794_ (.A(_02983_),
    .B(_02984_),
    .X(_02985_));
 sky130_fd_sc_hd__xor2_1 _22795_ (.A(_02136_),
    .B(_02985_),
    .X(_02986_));
 sky130_fd_sc_hd__xnor2_1 _22796_ (.A(_02978_),
    .B(_02986_),
    .Y(_02987_));
 sky130_fd_sc_hd__xnor2_1 _22797_ (.A(_02976_),
    .B(_02987_),
    .Y(_02988_));
 sky130_fd_sc_hd__nor2_1 _22798_ (.A(_02885_),
    .B(_02887_),
    .Y(_02989_));
 sky130_fd_sc_hd__and3_1 _22799_ (.A(_11237_),
    .B(_01547_),
    .C(_14570_),
    .X(_02990_));
 sky130_fd_sc_hd__o21ai_1 _22800_ (.A1(_11237_),
    .A2(_01547_),
    .B1(_14037_),
    .Y(_02991_));
 sky130_fd_sc_hd__nor2_1 _22801_ (.A(_02990_),
    .B(_02991_),
    .Y(_02992_));
 sky130_fd_sc_hd__o32a_1 _22802_ (.A1(_11137_),
    .A2(_02729_),
    .A3(_02866_),
    .B1(_02867_),
    .B2(_02732_),
    .X(_02993_));
 sky130_fd_sc_hd__xnor2_1 _22803_ (.A(_02992_),
    .B(_02993_),
    .Y(_02994_));
 sky130_fd_sc_hd__xnor2_1 _22804_ (.A(_02597_),
    .B(_02994_),
    .Y(_02995_));
 sky130_fd_sc_hd__or2b_1 _22805_ (.A(_02877_),
    .B_N(_02882_),
    .X(_02996_));
 sky130_fd_sc_hd__nand2_1 _22806_ (.A(_02876_),
    .B(_02883_),
    .Y(_02997_));
 sky130_fd_sc_hd__a31o_1 _22807_ (.A1(_11561_),
    .A2(_13817_),
    .A3(_02880_),
    .B1(_02879_),
    .X(_02998_));
 sky130_fd_sc_hd__o21ba_1 _22808_ (.A1(_02896_),
    .A2(_02899_),
    .B1_N(_02897_),
    .X(_02999_));
 sky130_fd_sc_hd__a22oi_1 _22809_ (.A1(_11925_),
    .A2(_13292_),
    .B1(_13605_),
    .B2(_11663_),
    .Y(_03000_));
 sky130_fd_sc_hd__and4_1 _22810_ (.A(_11555_),
    .B(_11658_),
    .C(\genblk1.pcpi_mul.rs1[29] ),
    .D(\genblk1.pcpi_mul.rs1[30] ),
    .X(_03001_));
 sky130_fd_sc_hd__nor2_1 _22811_ (.A(_03000_),
    .B(_03001_),
    .Y(_03002_));
 sky130_fd_sc_hd__nand2_1 _22812_ (.A(_11444_),
    .B(_14398_),
    .Y(_03003_));
 sky130_fd_sc_hd__xnor2_2 _22813_ (.A(_03002_),
    .B(_03003_),
    .Y(_03004_));
 sky130_fd_sc_hd__xnor2_1 _22814_ (.A(_02999_),
    .B(_03004_),
    .Y(_03005_));
 sky130_fd_sc_hd__xnor2_1 _22815_ (.A(_02998_),
    .B(_03005_),
    .Y(_03006_));
 sky130_fd_sc_hd__a21oi_1 _22816_ (.A1(_02996_),
    .A2(_02997_),
    .B1(_03006_),
    .Y(_03007_));
 sky130_fd_sc_hd__and3_1 _22817_ (.A(_02996_),
    .B(_02997_),
    .C(_03006_),
    .X(_03008_));
 sky130_fd_sc_hd__or3_1 _22818_ (.A(_02995_),
    .B(_03007_),
    .C(_03008_),
    .X(_03009_));
 sky130_fd_sc_hd__o21ai_1 _22819_ (.A1(_03007_),
    .A2(_03008_),
    .B1(_02995_),
    .Y(_03010_));
 sky130_fd_sc_hd__o211a_1 _22820_ (.A1(_02909_),
    .A2(_02911_),
    .B1(_03009_),
    .C1(_03010_),
    .X(_03011_));
 sky130_fd_sc_hd__a211o_1 _22821_ (.A1(_03009_),
    .A2(_03010_),
    .B1(_02909_),
    .C1(_02911_),
    .X(_03012_));
 sky130_fd_sc_hd__and2b_1 _22822_ (.A_N(_03011_),
    .B(_03012_),
    .X(_03013_));
 sky130_fd_sc_hd__xnor2_2 _22823_ (.A(_02989_),
    .B(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hd__or2b_1 _22824_ (.A(_02906_),
    .B_N(_02905_),
    .X(_03015_));
 sky130_fd_sc_hd__a21bo_2 _22825_ (.A1(_02900_),
    .A2(_02907_),
    .B1_N(_03015_),
    .X(_03016_));
 sky130_fd_sc_hd__or3_2 _22826_ (.A(_02914_),
    .B(_02917_),
    .C(_02918_),
    .X(_03017_));
 sky130_fd_sc_hd__a22oi_2 _22827_ (.A1(_01757_),
    .A2(_13286_),
    .B1(_01866_),
    .B2(_13936_),
    .Y(_03018_));
 sky130_fd_sc_hd__and4_1 _22828_ (.A(_01754_),
    .B(_01755_),
    .C(_13868_),
    .D(_01713_),
    .X(_03019_));
 sky130_fd_sc_hd__nor2_1 _22829_ (.A(_03018_),
    .B(_03019_),
    .Y(_03020_));
 sky130_fd_sc_hd__nand2_1 _22830_ (.A(_13711_),
    .B(_01717_),
    .Y(_03021_));
 sky130_fd_sc_hd__xnor2_1 _22831_ (.A(_03020_),
    .B(_03021_),
    .Y(_03022_));
 sky130_fd_sc_hd__a22oi_4 _22832_ (.A1(_14129_),
    .A2(_12830_),
    .B1(_13859_),
    .B2(_13942_),
    .Y(_03023_));
 sky130_fd_sc_hd__and4_1 _22833_ (.A(_12323_),
    .B(_13723_),
    .C(_12830_),
    .D(_12546_),
    .X(_03024_));
 sky130_fd_sc_hd__nor2_1 _22834_ (.A(_03023_),
    .B(_03024_),
    .Y(_03025_));
 sky130_fd_sc_hd__nand2_1 _22835_ (.A(_13720_),
    .B(_13861_),
    .Y(_03026_));
 sky130_fd_sc_hd__xnor2_1 _22836_ (.A(_03025_),
    .B(_03026_),
    .Y(_03027_));
 sky130_fd_sc_hd__o21ba_1 _22837_ (.A1(_02901_),
    .A2(_02904_),
    .B1_N(_02902_),
    .X(_03028_));
 sky130_fd_sc_hd__xnor2_1 _22838_ (.A(_03027_),
    .B(_03028_),
    .Y(_03029_));
 sky130_fd_sc_hd__xnor2_1 _22839_ (.A(_03022_),
    .B(_03029_),
    .Y(_03030_));
 sky130_fd_sc_hd__a21oi_1 _22840_ (.A1(_03017_),
    .A2(_02921_),
    .B1(_03030_),
    .Y(_03031_));
 sky130_fd_sc_hd__and3_1 _22841_ (.A(_03017_),
    .B(_02921_),
    .C(_03030_),
    .X(_03032_));
 sky130_fd_sc_hd__nor2_1 _22842_ (.A(_03031_),
    .B(_03032_),
    .Y(_03033_));
 sky130_fd_sc_hd__xor2_2 _22843_ (.A(_03016_),
    .B(_03033_),
    .X(_03034_));
 sky130_fd_sc_hd__o21ba_1 _22844_ (.A1(_02924_),
    .A2(_02927_),
    .B1_N(_02925_),
    .X(_03035_));
 sky130_fd_sc_hd__a22oi_2 _22845_ (.A1(_12271_),
    .A2(_13555_),
    .B1(_01601_),
    .B2(_12079_),
    .Y(_03036_));
 sky130_fd_sc_hd__and4_1 _22846_ (.A(_12144_),
    .B(_12273_),
    .C(_13558_),
    .D(_13740_),
    .X(_03037_));
 sky130_fd_sc_hd__nor2_1 _22847_ (.A(_03036_),
    .B(_03037_),
    .Y(_03038_));
 sky130_fd_sc_hd__nand2_1 _22848_ (.A(_13890_),
    .B(_14499_),
    .Y(_03039_));
 sky130_fd_sc_hd__xnor2_1 _22849_ (.A(_03038_),
    .B(_03039_),
    .Y(_03040_));
 sky130_fd_sc_hd__xnor2_2 _22850_ (.A(_03035_),
    .B(_03040_),
    .Y(_03041_));
 sky130_fd_sc_hd__o21ai_4 _22851_ (.A1(_02916_),
    .A2(_02918_),
    .B1(_03041_),
    .Y(_03042_));
 sky130_fd_sc_hd__or3_1 _22852_ (.A(_02916_),
    .B(_02918_),
    .C(_03041_),
    .X(_03043_));
 sky130_fd_sc_hd__and2_2 _22853_ (.A(_03042_),
    .B(_03043_),
    .X(_03044_));
 sky130_fd_sc_hd__a22oi_2 _22854_ (.A1(_11950_),
    .A2(_13970_),
    .B1(_13972_),
    .B2(_11820_),
    .Y(_03045_));
 sky130_fd_sc_hd__and4_1 _22855_ (.A(_13918_),
    .B(_13679_),
    .C(_13764_),
    .D(_13765_),
    .X(_03046_));
 sky130_fd_sc_hd__nor2_1 _22856_ (.A(_03045_),
    .B(_03046_),
    .Y(_03047_));
 sky130_fd_sc_hd__nand2_1 _22857_ (.A(_14457_),
    .B(_13056_),
    .Y(_03048_));
 sky130_fd_sc_hd__xnor2_2 _22858_ (.A(_03047_),
    .B(_03048_),
    .Y(_03049_));
 sky130_fd_sc_hd__and2b_1 _22859_ (.A_N(_11481_),
    .B(_02237_),
    .X(_03050_));
 sky130_fd_sc_hd__nand2_1 _22860_ (.A(_11489_),
    .B(_14167_),
    .Y(_03051_));
 sky130_fd_sc_hd__xnor2_2 _22861_ (.A(_03050_),
    .B(_03051_),
    .Y(_03052_));
 sky130_fd_sc_hd__nand2_1 _22862_ (.A(_13695_),
    .B(_14342_),
    .Y(_03053_));
 sky130_fd_sc_hd__xnor2_2 _22863_ (.A(_03052_),
    .B(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__and3_1 _22864_ (.A(_12561_),
    .B(_01620_),
    .C(_02930_),
    .X(_03055_));
 sky130_fd_sc_hd__a31o_1 _22865_ (.A1(_11826_),
    .A2(_13752_),
    .A3(_02932_),
    .B1(_03055_),
    .X(_03056_));
 sky130_fd_sc_hd__xor2_2 _22866_ (.A(_03054_),
    .B(_03056_),
    .X(_03057_));
 sky130_fd_sc_hd__xnor2_2 _22867_ (.A(_03049_),
    .B(_03057_),
    .Y(_03058_));
 sky130_fd_sc_hd__nand2_1 _22868_ (.A(_02933_),
    .B(_02935_),
    .Y(_03059_));
 sky130_fd_sc_hd__a21boi_2 _22869_ (.A1(_02928_),
    .A2(_02936_),
    .B1_N(_03059_),
    .Y(_03060_));
 sky130_fd_sc_hd__xnor2_2 _22870_ (.A(_03058_),
    .B(_03060_),
    .Y(_03061_));
 sky130_fd_sc_hd__xnor2_4 _22871_ (.A(_03044_),
    .B(_03061_),
    .Y(_03062_));
 sky130_fd_sc_hd__nand2_1 _22872_ (.A(_02937_),
    .B(_02939_),
    .Y(_03063_));
 sky130_fd_sc_hd__nor2_1 _22873_ (.A(_02937_),
    .B(_02939_),
    .Y(_03064_));
 sky130_fd_sc_hd__a21oi_4 _22874_ (.A1(_02923_),
    .A2(_03063_),
    .B1(_03064_),
    .Y(_03065_));
 sky130_fd_sc_hd__xnor2_2 _22875_ (.A(_03062_),
    .B(_03065_),
    .Y(_03066_));
 sky130_fd_sc_hd__xnor2_2 _22876_ (.A(_03034_),
    .B(_03066_),
    .Y(_03067_));
 sky130_fd_sc_hd__and2b_1 _22877_ (.A_N(_02944_),
    .B(_02941_),
    .X(_03068_));
 sky130_fd_sc_hd__a21oi_4 _22878_ (.A1(_02913_),
    .A2(_02945_),
    .B1(_03068_),
    .Y(_03069_));
 sky130_fd_sc_hd__xor2_2 _22879_ (.A(_03067_),
    .B(_03069_),
    .X(_03070_));
 sky130_fd_sc_hd__xor2_2 _22880_ (.A(_03014_),
    .B(_03070_),
    .X(_03071_));
 sky130_fd_sc_hd__nor2_1 _22881_ (.A(_02946_),
    .B(_02948_),
    .Y(_03072_));
 sky130_fd_sc_hd__a21o_1 _22882_ (.A1(_02892_),
    .A2(_02949_),
    .B1(_03072_),
    .X(_03073_));
 sky130_fd_sc_hd__xor2_1 _22883_ (.A(_03071_),
    .B(_03073_),
    .X(_03074_));
 sky130_fd_sc_hd__xnor2_1 _22884_ (.A(_02988_),
    .B(_03074_),
    .Y(_03075_));
 sky130_fd_sc_hd__and2b_1 _22885_ (.A_N(_02952_),
    .B(_02950_),
    .X(_03076_));
 sky130_fd_sc_hd__a21o_1 _22886_ (.A1(_02862_),
    .A2(_02953_),
    .B1(_03076_),
    .X(_03077_));
 sky130_fd_sc_hd__xor2_1 _22887_ (.A(_03075_),
    .B(_03077_),
    .X(_03078_));
 sky130_fd_sc_hd__xnor2_2 _22888_ (.A(_02974_),
    .B(_03078_),
    .Y(_03079_));
 sky130_fd_sc_hd__nor2_1 _22889_ (.A(_02954_),
    .B(_02956_),
    .Y(_03080_));
 sky130_fd_sc_hd__nand2_1 _22890_ (.A(_02954_),
    .B(_02956_),
    .Y(_03081_));
 sky130_fd_sc_hd__o21a_1 _22891_ (.A1(_02842_),
    .A2(_03080_),
    .B1(_03081_),
    .X(_03082_));
 sky130_fd_sc_hd__xnor2_2 _22892_ (.A(_03079_),
    .B(_03082_),
    .Y(_03083_));
 sky130_fd_sc_hd__xnor2_4 _22893_ (.A(_02970_),
    .B(_03083_),
    .Y(_03084_));
 sky130_fd_sc_hd__and2b_1 _22894_ (.A_N(_02961_),
    .B(_02958_),
    .X(_03085_));
 sky130_fd_sc_hd__a21oi_2 _22895_ (.A1(_02838_),
    .A2(_02962_),
    .B1(_03085_),
    .Y(_03086_));
 sky130_fd_sc_hd__xor2_4 _22896_ (.A(_03084_),
    .B(_03086_),
    .X(_03087_));
 sky130_fd_sc_hd__or3b_1 _22897_ (.A(_02966_),
    .B(_02830_),
    .C_N(_02964_),
    .X(_03088_));
 sky130_fd_sc_hd__a21o_1 _22898_ (.A1(_02968_),
    .A2(_02964_),
    .B1(_02966_),
    .X(_03089_));
 sky130_fd_sc_hd__o21a_2 _22899_ (.A1(_02835_),
    .A2(_03088_),
    .B1(_03089_),
    .X(_03090_));
 sky130_fd_sc_hd__xnor2_4 _22900_ (.A(_03087_),
    .B(_03090_),
    .Y(_00092_));
 sky130_fd_sc_hd__or2b_1 _22901_ (.A(_03082_),
    .B_N(_03079_),
    .X(_03091_));
 sky130_fd_sc_hd__nand2_1 _22902_ (.A(_02970_),
    .B(_03083_),
    .Y(_03092_));
 sky130_fd_sc_hd__a21oi_1 _22903_ (.A1(_02971_),
    .A2(_02972_),
    .B1(_02567_),
    .Y(_03093_));
 sky130_fd_sc_hd__or2b_1 _22904_ (.A(_02978_),
    .B_N(_02986_),
    .X(_03094_));
 sky130_fd_sc_hd__nand2_1 _22905_ (.A(_02976_),
    .B(_02987_),
    .Y(_03095_));
 sky130_fd_sc_hd__a21oi_1 _22906_ (.A1(_03094_),
    .A2(_03095_),
    .B1(_02287_),
    .Y(_03096_));
 sky130_fd_sc_hd__and3_1 _22907_ (.A(_02132_),
    .B(_03094_),
    .C(_03095_),
    .X(_03097_));
 sky130_fd_sc_hd__or2_1 _22908_ (.A(_03096_),
    .B(_03097_),
    .X(_03098_));
 sky130_fd_sc_hd__or2b_1 _22909_ (.A(_02984_),
    .B_N(_02983_),
    .X(_03099_));
 sky130_fd_sc_hd__o21ai_1 _22910_ (.A1(_02433_),
    .A2(_02985_),
    .B1(_03099_),
    .Y(_03100_));
 sky130_fd_sc_hd__or3b_1 _22911_ (.A(_02989_),
    .B(_03011_),
    .C_N(_03012_),
    .X(_03101_));
 sky130_fd_sc_hd__or2b_1 _22912_ (.A(_03011_),
    .B_N(_03101_),
    .X(_03102_));
 sky130_fd_sc_hd__o21ai_1 _22913_ (.A1(_02854_),
    .A2(_02982_),
    .B1(_02980_),
    .Y(_03103_));
 sky130_fd_sc_hd__and2_1 _22914_ (.A(_11137_),
    .B(_02990_),
    .X(_03104_));
 sky130_fd_sc_hd__a21oi_1 _22915_ (.A1(_02598_),
    .A2(_02994_),
    .B1(_03104_),
    .Y(_03105_));
 sky130_fd_sc_hd__nor2_1 _22916_ (.A(_02848_),
    .B(_02854_),
    .Y(_03106_));
 sky130_fd_sc_hd__or2_1 _22917_ (.A(_02445_),
    .B(_02852_),
    .X(_03107_));
 sky130_fd_sc_hd__or2b_1 _22918_ (.A(_03106_),
    .B_N(_03107_),
    .X(_03108_));
 sky130_fd_sc_hd__xnor2_1 _22919_ (.A(_03105_),
    .B(_03108_),
    .Y(_03109_));
 sky130_fd_sc_hd__xnor2_1 _22920_ (.A(_03103_),
    .B(_03109_),
    .Y(_03110_));
 sky130_fd_sc_hd__xnor2_1 _22921_ (.A(_02137_),
    .B(_03110_),
    .Y(_03111_));
 sky130_fd_sc_hd__xnor2_1 _22922_ (.A(_03102_),
    .B(_03111_),
    .Y(_03112_));
 sky130_fd_sc_hd__xor2_1 _22923_ (.A(_03100_),
    .B(_03112_),
    .X(_03113_));
 sky130_fd_sc_hd__or2b_1 _22924_ (.A(_03007_),
    .B_N(_03009_),
    .X(_03114_));
 sky130_fd_sc_hd__a21o_1 _22925_ (.A1(_03016_),
    .A2(_03033_),
    .B1(_03031_),
    .X(_03115_));
 sky130_fd_sc_hd__nand2_1 _22926_ (.A(_02732_),
    .B(_02991_),
    .Y(_03116_));
 sky130_fd_sc_hd__nand2b_4 _22927_ (.A_N(_03104_),
    .B(_03116_),
    .Y(_03117_));
 sky130_fd_sc_hd__xor2_4 _22928_ (.A(_02598_),
    .B(_03117_),
    .X(_03118_));
 sky130_fd_sc_hd__or2b_1 _22929_ (.A(_02999_),
    .B_N(_03004_),
    .X(_03119_));
 sky130_fd_sc_hd__nand2_1 _22930_ (.A(_02998_),
    .B(_03005_),
    .Y(_03120_));
 sky130_fd_sc_hd__a31o_1 _22931_ (.A1(_14099_),
    .A2(_14212_),
    .A3(_03002_),
    .B1(_03001_),
    .X(_03121_));
 sky130_fd_sc_hd__o21ba_1 _22932_ (.A1(_03018_),
    .A2(_03021_),
    .B1_N(_03019_),
    .X(_03122_));
 sky130_fd_sc_hd__a22oi_4 _22933_ (.A1(_11782_),
    .A2(_13606_),
    .B1(_14398_),
    .B2(_11664_),
    .Y(_03123_));
 sky130_fd_sc_hd__and4_1 _22934_ (.A(_11556_),
    .B(_11665_),
    .C(_13605_),
    .D(\genblk1.pcpi_mul.rs1[31] ),
    .X(_03124_));
 sky130_fd_sc_hd__nor2_1 _22935_ (.A(_03123_),
    .B(_03124_),
    .Y(_03125_));
 sky130_fd_sc_hd__nand2_2 _22936_ (.A(_11560_),
    .B(_14026_),
    .Y(_03126_));
 sky130_fd_sc_hd__xnor2_1 _22937_ (.A(_03125_),
    .B(_03126_),
    .Y(_03127_));
 sky130_fd_sc_hd__xnor2_1 _22938_ (.A(_03122_),
    .B(_03127_),
    .Y(_03128_));
 sky130_fd_sc_hd__xnor2_1 _22939_ (.A(_03121_),
    .B(_03128_),
    .Y(_03129_));
 sky130_fd_sc_hd__a21oi_1 _22940_ (.A1(_03119_),
    .A2(_03120_),
    .B1(_03129_),
    .Y(_03130_));
 sky130_fd_sc_hd__and3_1 _22941_ (.A(_03119_),
    .B(_03120_),
    .C(_03129_),
    .X(_03131_));
 sky130_fd_sc_hd__or2_1 _22942_ (.A(_03130_),
    .B(_03131_),
    .X(_03132_));
 sky130_fd_sc_hd__xnor2_1 _22943_ (.A(_03118_),
    .B(_03132_),
    .Y(_03133_));
 sky130_fd_sc_hd__xor2_1 _22944_ (.A(_03115_),
    .B(_03133_),
    .X(_03134_));
 sky130_fd_sc_hd__xnor2_2 _22945_ (.A(_03114_),
    .B(_03134_),
    .Y(_03135_));
 sky130_fd_sc_hd__and2b_1 _22946_ (.A_N(_03028_),
    .B(_03027_),
    .X(_03136_));
 sky130_fd_sc_hd__and2_1 _22947_ (.A(_03022_),
    .B(_03029_),
    .X(_03137_));
 sky130_fd_sc_hd__or2b_2 _22948_ (.A(_03035_),
    .B_N(_03040_),
    .X(_03138_));
 sky130_fd_sc_hd__a22oi_2 _22949_ (.A1(_01583_),
    .A2(_14059_),
    .B1(_01844_),
    .B2(_11892_),
    .Y(_03139_));
 sky130_fd_sc_hd__and4_1 _22950_ (.A(_01582_),
    .B(_01757_),
    .C(_01866_),
    .D(_13612_),
    .X(_03140_));
 sky130_fd_sc_hd__nor2_1 _22951_ (.A(_03139_),
    .B(_03140_),
    .Y(_03141_));
 sky130_fd_sc_hd__nand2_1 _22952_ (.A(_11772_),
    .B(_13815_),
    .Y(_03142_));
 sky130_fd_sc_hd__xnor2_1 _22953_ (.A(_03141_),
    .B(_03142_),
    .Y(_03143_));
 sky130_fd_sc_hd__a22oi_2 _22954_ (.A1(_14310_),
    .A2(_14076_),
    .B1(_13864_),
    .B2(_14132_),
    .Y(_03144_));
 sky130_fd_sc_hd__and4_1 _22955_ (.A(_13942_),
    .B(_13721_),
    .C(_13859_),
    .D(_13637_),
    .X(_03145_));
 sky130_fd_sc_hd__nor2_1 _22956_ (.A(_03144_),
    .B(_03145_),
    .Y(_03146_));
 sky130_fd_sc_hd__nand2_1 _22957_ (.A(_13720_),
    .B(_14438_),
    .Y(_03147_));
 sky130_fd_sc_hd__xnor2_1 _22958_ (.A(_03146_),
    .B(_03147_),
    .Y(_03148_));
 sky130_fd_sc_hd__o21ba_1 _22959_ (.A1(_03023_),
    .A2(_03026_),
    .B1_N(_03024_),
    .X(_03149_));
 sky130_fd_sc_hd__xnor2_1 _22960_ (.A(_03148_),
    .B(_03149_),
    .Y(_03150_));
 sky130_fd_sc_hd__xnor2_1 _22961_ (.A(_03143_),
    .B(_03150_),
    .Y(_03151_));
 sky130_fd_sc_hd__a21o_1 _22962_ (.A1(_03138_),
    .A2(_03042_),
    .B1(_03151_),
    .X(_03152_));
 sky130_fd_sc_hd__nand3_1 _22963_ (.A(_03138_),
    .B(_03042_),
    .C(_03151_),
    .Y(_03153_));
 sky130_fd_sc_hd__o211ai_2 _22964_ (.A1(_03136_),
    .A2(_03137_),
    .B1(_03152_),
    .C1(_03153_),
    .Y(_03154_));
 sky130_fd_sc_hd__a211o_1 _22965_ (.A1(_03152_),
    .A2(_03153_),
    .B1(_03136_),
    .C1(_03137_),
    .X(_03155_));
 sky130_fd_sc_hd__and2_1 _22966_ (.A(_03154_),
    .B(_03155_),
    .X(_03156_));
 sky130_fd_sc_hd__o21ba_2 _22967_ (.A1(_03036_),
    .A2(_03039_),
    .B1_N(_03037_),
    .X(_03157_));
 sky130_fd_sc_hd__o21ba_2 _22968_ (.A1(_03045_),
    .A2(_03048_),
    .B1_N(_03046_),
    .X(_03158_));
 sky130_fd_sc_hd__clkbuf_2 _22969_ (.A(_13744_),
    .X(_03159_));
 sky130_fd_sc_hd__a22oi_1 _22970_ (.A1(_14269_),
    .A2(_12772_),
    .B1(_03159_),
    .B2(_13668_),
    .Y(_03160_));
 sky130_fd_sc_hd__and4_1 _22971_ (.A(_12543_),
    .B(_12694_),
    .C(_13739_),
    .D(_13741_),
    .X(_03161_));
 sky130_fd_sc_hd__nor2_1 _22972_ (.A(_03160_),
    .B(_03161_),
    .Y(_03162_));
 sky130_fd_sc_hd__nand2_1 _22973_ (.A(_13888_),
    .B(_12586_),
    .Y(_03163_));
 sky130_fd_sc_hd__xnor2_1 _22974_ (.A(_03162_),
    .B(_03163_),
    .Y(_03164_));
 sky130_fd_sc_hd__xnor2_1 _22975_ (.A(_03158_),
    .B(_03164_),
    .Y(_03165_));
 sky130_fd_sc_hd__xnor2_2 _22976_ (.A(_03157_),
    .B(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hd__and2b_2 _22977_ (.A_N(_11961_),
    .B(_01618_),
    .X(_03167_));
 sky130_fd_sc_hd__nand2_2 _22978_ (.A(_11699_),
    .B(_01620_),
    .Y(_03168_));
 sky130_fd_sc_hd__xnor2_4 _22979_ (.A(_03167_),
    .B(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__nand2_2 _22980_ (.A(_12075_),
    .B(_14343_),
    .Y(_03170_));
 sky130_fd_sc_hd__xnor2_4 _22981_ (.A(_03169_),
    .B(_03170_),
    .Y(_03171_));
 sky130_fd_sc_hd__and3_1 _22982_ (.A(_11491_),
    .B(_01625_),
    .C(_03050_),
    .X(_03172_));
 sky130_fd_sc_hd__a31o_2 _22983_ (.A1(_11954_),
    .A2(_01624_),
    .A3(_03052_),
    .B1(_03172_),
    .X(_03173_));
 sky130_fd_sc_hd__xor2_2 _22984_ (.A(_03171_),
    .B(_03173_),
    .X(_03174_));
 sky130_fd_sc_hd__clkbuf_2 _22985_ (.A(_13972_),
    .X(_03175_));
 sky130_fd_sc_hd__a22oi_2 _22986_ (.A1(_12278_),
    .A2(_13229_),
    .B1(_03175_),
    .B2(_14283_),
    .Y(_03176_));
 sky130_fd_sc_hd__and4_1 _22987_ (.A(_13904_),
    .B(_12278_),
    .C(_13224_),
    .D(_14510_),
    .X(_03177_));
 sky130_fd_sc_hd__nor2_2 _22988_ (.A(_03176_),
    .B(_03177_),
    .Y(_03178_));
 sky130_fd_sc_hd__clkbuf_2 _22989_ (.A(_13056_),
    .X(_03179_));
 sky130_fd_sc_hd__nand2_2 _22990_ (.A(_01558_),
    .B(_03179_),
    .Y(_03180_));
 sky130_fd_sc_hd__xnor2_4 _22991_ (.A(_03178_),
    .B(_03180_),
    .Y(_03181_));
 sky130_fd_sc_hd__xnor2_2 _22992_ (.A(_03174_),
    .B(_03181_),
    .Y(_03182_));
 sky130_fd_sc_hd__and2_1 _22993_ (.A(_03054_),
    .B(_03056_),
    .X(_03183_));
 sky130_fd_sc_hd__a21o_2 _22994_ (.A1(_03049_),
    .A2(_03057_),
    .B1(_03183_),
    .X(_03184_));
 sky130_fd_sc_hd__xnor2_2 _22995_ (.A(_03182_),
    .B(_03184_),
    .Y(_03185_));
 sky130_fd_sc_hd__xor2_2 _22996_ (.A(_03166_),
    .B(_03185_),
    .X(_03186_));
 sky130_fd_sc_hd__nand2_1 _22997_ (.A(_03058_),
    .B(_03060_),
    .Y(_03187_));
 sky130_fd_sc_hd__nor2_1 _22998_ (.A(_03058_),
    .B(_03060_),
    .Y(_03188_));
 sky130_fd_sc_hd__a21oi_4 _22999_ (.A1(_03044_),
    .A2(_03187_),
    .B1(_03188_),
    .Y(_03189_));
 sky130_fd_sc_hd__xnor2_2 _23000_ (.A(_03186_),
    .B(_03189_),
    .Y(_03190_));
 sky130_fd_sc_hd__xnor2_2 _23001_ (.A(_03156_),
    .B(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__and2b_1 _23002_ (.A_N(_03065_),
    .B(_03062_),
    .X(_03192_));
 sky130_fd_sc_hd__a21oi_2 _23003_ (.A1(_03034_),
    .A2(_03066_),
    .B1(_03192_),
    .Y(_03193_));
 sky130_fd_sc_hd__xnor2_1 _23004_ (.A(_03191_),
    .B(_03193_),
    .Y(_03194_));
 sky130_fd_sc_hd__xor2_2 _23005_ (.A(_03135_),
    .B(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__nor2_1 _23006_ (.A(_03067_),
    .B(_03069_),
    .Y(_03196_));
 sky130_fd_sc_hd__a21oi_1 _23007_ (.A1(_03014_),
    .A2(_03070_),
    .B1(_03196_),
    .Y(_03197_));
 sky130_fd_sc_hd__xnor2_1 _23008_ (.A(_03195_),
    .B(_03197_),
    .Y(_03198_));
 sky130_fd_sc_hd__xnor2_1 _23009_ (.A(_03113_),
    .B(_03198_),
    .Y(_03199_));
 sky130_fd_sc_hd__nor2_1 _23010_ (.A(_03071_),
    .B(_03073_),
    .Y(_03200_));
 sky130_fd_sc_hd__nand2_1 _23011_ (.A(_03071_),
    .B(_03073_),
    .Y(_03201_));
 sky130_fd_sc_hd__o21a_1 _23012_ (.A1(_02988_),
    .A2(_03200_),
    .B1(_03201_),
    .X(_03202_));
 sky130_fd_sc_hd__xor2_1 _23013_ (.A(_03199_),
    .B(_03202_),
    .X(_03203_));
 sky130_fd_sc_hd__xnor2_1 _23014_ (.A(_03098_),
    .B(_03203_),
    .Y(_03204_));
 sky130_fd_sc_hd__nor2_1 _23015_ (.A(_03075_),
    .B(_03077_),
    .Y(_03205_));
 sky130_fd_sc_hd__nand2_1 _23016_ (.A(_03075_),
    .B(_03077_),
    .Y(_03206_));
 sky130_fd_sc_hd__o21ai_1 _23017_ (.A1(_02974_),
    .A2(_03205_),
    .B1(_03206_),
    .Y(_03207_));
 sky130_fd_sc_hd__xor2_1 _23018_ (.A(_03204_),
    .B(_03207_),
    .X(_03208_));
 sky130_fd_sc_hd__xnor2_1 _23019_ (.A(_03093_),
    .B(_03208_),
    .Y(_03209_));
 sky130_fd_sc_hd__nand3_1 _23020_ (.A(_03091_),
    .B(_03092_),
    .C(_03209_),
    .Y(_03210_));
 sky130_vsdinv _23021_ (.A(_03210_),
    .Y(_03211_));
 sky130_fd_sc_hd__a21oi_2 _23022_ (.A1(_03091_),
    .A2(_03092_),
    .B1(_03209_),
    .Y(_03212_));
 sky130_fd_sc_hd__nor2_2 _23023_ (.A(_03211_),
    .B(_03212_),
    .Y(_03213_));
 sky130_fd_sc_hd__nor2_1 _23024_ (.A(_03084_),
    .B(_03086_),
    .Y(_03214_));
 sky130_fd_sc_hd__and2b_1 _23025_ (.A_N(_03090_),
    .B(_03087_),
    .X(_03215_));
 sky130_fd_sc_hd__nor2_2 _23026_ (.A(_03214_),
    .B(_03215_),
    .Y(_03216_));
 sky130_fd_sc_hd__xnor2_4 _23027_ (.A(_03213_),
    .B(_03216_),
    .Y(_00093_));
 sky130_fd_sc_hd__nand2_1 _23028_ (.A(_03102_),
    .B(_03111_),
    .Y(_03217_));
 sky130_fd_sc_hd__or2b_1 _23029_ (.A(_03112_),
    .B_N(_03100_),
    .X(_03218_));
 sky130_fd_sc_hd__clkbuf_2 _23030_ (.A(_02425_),
    .X(_03219_));
 sky130_fd_sc_hd__a21oi_1 _23031_ (.A1(_03217_),
    .A2(_03218_),
    .B1(_03219_),
    .Y(_03220_));
 sky130_fd_sc_hd__and3_1 _23032_ (.A(_02426_),
    .B(_03217_),
    .C(_03218_),
    .X(_03221_));
 sky130_fd_sc_hd__or2_1 _23033_ (.A(_03220_),
    .B(_03221_),
    .X(_03222_));
 sky130_fd_sc_hd__or2_1 _23034_ (.A(_02854_),
    .B(_02982_),
    .X(_03223_));
 sky130_fd_sc_hd__a21oi_1 _23035_ (.A1(_02980_),
    .A2(_03223_),
    .B1(_03109_),
    .Y(_03224_));
 sky130_fd_sc_hd__or2b_1 _23036_ (.A(_02433_),
    .B_N(_03110_),
    .X(_03225_));
 sky130_fd_sc_hd__or2b_1 _23037_ (.A(_03224_),
    .B_N(_03225_),
    .X(_03226_));
 sky130_fd_sc_hd__and2b_1 _23038_ (.A_N(_03133_),
    .B(_03115_),
    .X(_03227_));
 sky130_fd_sc_hd__and2b_1 _23039_ (.A_N(_03134_),
    .B(_03114_),
    .X(_03228_));
 sky130_fd_sc_hd__a21o_1 _23040_ (.A1(_02598_),
    .A2(_03116_),
    .B1(_03104_),
    .X(_03229_));
 sky130_fd_sc_hd__or2_1 _23041_ (.A(_03105_),
    .B(_03106_),
    .X(_03230_));
 sky130_fd_sc_hd__nor2_1 _23042_ (.A(_03107_),
    .B(_03229_),
    .Y(_03231_));
 sky130_fd_sc_hd__a31o_1 _23043_ (.A1(_03107_),
    .A2(_03229_),
    .A3(_03230_),
    .B1(_03231_),
    .X(_03232_));
 sky130_fd_sc_hd__xor2_1 _23044_ (.A(_02137_),
    .B(_03232_),
    .X(_03233_));
 sky130_fd_sc_hd__o21ai_1 _23045_ (.A1(_03227_),
    .A2(_03228_),
    .B1(_03233_),
    .Y(_03234_));
 sky130_fd_sc_hd__or3_1 _23046_ (.A(_03227_),
    .B(_03228_),
    .C(_03233_),
    .X(_03235_));
 sky130_fd_sc_hd__and2_1 _23047_ (.A(_03234_),
    .B(_03235_),
    .X(_03236_));
 sky130_fd_sc_hd__xnor2_1 _23048_ (.A(_03226_),
    .B(_03236_),
    .Y(_03237_));
 sky130_fd_sc_hd__clkbuf_2 _23049_ (.A(_03118_),
    .X(_03238_));
 sky130_fd_sc_hd__o21ba_1 _23050_ (.A1(_03238_),
    .A2(_03132_),
    .B1_N(_03130_),
    .X(_03239_));
 sky130_fd_sc_hd__xnor2_4 _23051_ (.A(_02598_),
    .B(_03117_),
    .Y(_03240_));
 sky130_fd_sc_hd__or2b_1 _23052_ (.A(_03122_),
    .B_N(_03127_),
    .X(_03241_));
 sky130_fd_sc_hd__nand2_1 _23053_ (.A(_03121_),
    .B(_03128_),
    .Y(_03242_));
 sky130_fd_sc_hd__o21ba_1 _23054_ (.A1(_03139_),
    .A2(_03142_),
    .B1_N(_03140_),
    .X(_03243_));
 sky130_vsdinv _23055_ (.A(_03126_),
    .Y(_03244_));
 sky130_fd_sc_hd__and3_2 _23056_ (.A(_11556_),
    .B(_11665_),
    .C(_14024_),
    .X(_03245_));
 sky130_fd_sc_hd__a22o_1 _23057_ (.A1(_11666_),
    .A2(_13830_),
    .B1(_14026_),
    .B2(_11557_),
    .X(_03246_));
 sky130_fd_sc_hd__a21bo_1 _23058_ (.A1(_14211_),
    .A2(_03245_),
    .B1_N(_03246_),
    .X(_03247_));
 sky130_fd_sc_hd__xnor2_1 _23059_ (.A(_03244_),
    .B(_03247_),
    .Y(_03248_));
 sky130_fd_sc_hd__xnor2_1 _23060_ (.A(_03243_),
    .B(_03248_),
    .Y(_03249_));
 sky130_fd_sc_hd__a21oi_1 _23061_ (.A1(_03125_),
    .A2(_03244_),
    .B1(_03124_),
    .Y(_03250_));
 sky130_fd_sc_hd__xor2_1 _23062_ (.A(_03249_),
    .B(_03250_),
    .X(_03251_));
 sky130_fd_sc_hd__a21oi_1 _23063_ (.A1(_03241_),
    .A2(_03242_),
    .B1(_03251_),
    .Y(_03252_));
 sky130_fd_sc_hd__and3_1 _23064_ (.A(_03241_),
    .B(_03242_),
    .C(_03251_),
    .X(_03253_));
 sky130_fd_sc_hd__nor2_1 _23065_ (.A(_03252_),
    .B(_03253_),
    .Y(_03254_));
 sky130_fd_sc_hd__xnor2_1 _23066_ (.A(_03240_),
    .B(_03254_),
    .Y(_03255_));
 sky130_fd_sc_hd__a21oi_1 _23067_ (.A1(_03152_),
    .A2(_03154_),
    .B1(_03255_),
    .Y(_03256_));
 sky130_fd_sc_hd__and3_1 _23068_ (.A(_03152_),
    .B(_03154_),
    .C(_03255_),
    .X(_03257_));
 sky130_fd_sc_hd__nor2_1 _23069_ (.A(_03256_),
    .B(_03257_),
    .Y(_03258_));
 sky130_fd_sc_hd__xor2_1 _23070_ (.A(_03239_),
    .B(_03258_),
    .X(_03259_));
 sky130_fd_sc_hd__or2b_1 _23071_ (.A(_03149_),
    .B_N(_03148_),
    .X(_03260_));
 sky130_fd_sc_hd__a21bo_1 _23072_ (.A1(_03143_),
    .A2(_03150_),
    .B1_N(_03260_),
    .X(_03261_));
 sky130_fd_sc_hd__or2b_1 _23073_ (.A(_03158_),
    .B_N(_03164_),
    .X(_03262_));
 sky130_fd_sc_hd__or2b_1 _23074_ (.A(_03157_),
    .B_N(_03165_),
    .X(_03263_));
 sky130_fd_sc_hd__a22oi_1 _23075_ (.A1(_01757_),
    .A2(_13612_),
    .B1(_01870_),
    .B2(_01582_),
    .Y(_03264_));
 sky130_fd_sc_hd__and4_1 _23076_ (.A(_01754_),
    .B(_01755_),
    .C(_01516_),
    .D(_14033_),
    .X(_03265_));
 sky130_fd_sc_hd__nor2_1 _23077_ (.A(_03264_),
    .B(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__nand2_1 _23078_ (.A(_11773_),
    .B(_14023_),
    .Y(_03267_));
 sky130_fd_sc_hd__xnor2_1 _23079_ (.A(_03266_),
    .B(_03267_),
    .Y(_03268_));
 sky130_fd_sc_hd__a22oi_2 _23080_ (.A1(_13945_),
    .A2(_13864_),
    .B1(_13286_),
    .B2(_12324_),
    .Y(_03269_));
 sky130_fd_sc_hd__and4_1 _23081_ (.A(_14132_),
    .B(_14310_),
    .C(_13637_),
    .D(_14056_),
    .X(_03270_));
 sky130_fd_sc_hd__nor2_1 _23082_ (.A(_03269_),
    .B(_03270_),
    .Y(_03271_));
 sky130_fd_sc_hd__nand2_1 _23083_ (.A(_12228_),
    .B(_14059_),
    .Y(_03272_));
 sky130_fd_sc_hd__xnor2_1 _23084_ (.A(_03271_),
    .B(_03272_),
    .Y(_03273_));
 sky130_fd_sc_hd__o21ba_1 _23085_ (.A1(_03144_),
    .A2(_03147_),
    .B1_N(_03145_),
    .X(_03274_));
 sky130_fd_sc_hd__xnor2_1 _23086_ (.A(_03273_),
    .B(_03274_),
    .Y(_03275_));
 sky130_fd_sc_hd__xnor2_1 _23087_ (.A(_03268_),
    .B(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__a21oi_1 _23088_ (.A1(_03262_),
    .A2(_03263_),
    .B1(_03276_),
    .Y(_03277_));
 sky130_fd_sc_hd__and3_1 _23089_ (.A(_03262_),
    .B(_03263_),
    .C(_03276_),
    .X(_03278_));
 sky130_fd_sc_hd__or2_1 _23090_ (.A(_03277_),
    .B(_03278_),
    .X(_03279_));
 sky130_fd_sc_hd__xnor2_1 _23091_ (.A(_03261_),
    .B(_03279_),
    .Y(_03280_));
 sky130_fd_sc_hd__and2b_1 _23092_ (.A_N(_11699_),
    .B(_13803_),
    .X(_03281_));
 sky130_fd_sc_hd__nand2_1 _23093_ (.A(_11820_),
    .B(_13757_),
    .Y(_03282_));
 sky130_fd_sc_hd__xnor2_2 _23094_ (.A(_03281_),
    .B(_03282_),
    .Y(_03283_));
 sky130_fd_sc_hd__nand2_1 _23095_ (.A(_14283_),
    .B(_01624_),
    .Y(_03284_));
 sky130_fd_sc_hd__xnor2_2 _23096_ (.A(_03283_),
    .B(_03284_),
    .Y(_03285_));
 sky130_fd_sc_hd__buf_2 _23097_ (.A(_13752_),
    .X(_03286_));
 sky130_fd_sc_hd__clkbuf_2 _23098_ (.A(_13757_),
    .X(_03287_));
 sky130_fd_sc_hd__and3_1 _23099_ (.A(_11954_),
    .B(_03287_),
    .C(_03167_),
    .X(_03288_));
 sky130_fd_sc_hd__a31o_2 _23100_ (.A1(_13919_),
    .A2(_03286_),
    .A3(_03169_),
    .B1(_03288_),
    .X(_03289_));
 sky130_fd_sc_hd__xor2_2 _23101_ (.A(_03285_),
    .B(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__a22oi_1 _23102_ (.A1(_13667_),
    .A2(_13229_),
    .B1(_01613_),
    .B2(_12278_),
    .Y(_03291_));
 sky130_fd_sc_hd__and4_1 _23103_ (.A(_13674_),
    .B(_12413_),
    .C(_13224_),
    .D(_13972_),
    .X(_03292_));
 sky130_fd_sc_hd__nor2_1 _23104_ (.A(_03291_),
    .B(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hd__nand2_1 _23105_ (.A(_13893_),
    .B(_13056_),
    .Y(_03294_));
 sky130_fd_sc_hd__xnor2_2 _23106_ (.A(_03293_),
    .B(_03294_),
    .Y(_03295_));
 sky130_fd_sc_hd__xnor2_2 _23107_ (.A(_03290_),
    .B(_03295_),
    .Y(_03296_));
 sky130_fd_sc_hd__and2_1 _23108_ (.A(_03171_),
    .B(_03173_),
    .X(_03297_));
 sky130_fd_sc_hd__a21o_1 _23109_ (.A1(_03174_),
    .A2(_03181_),
    .B1(_03297_),
    .X(_03298_));
 sky130_fd_sc_hd__xnor2_1 _23110_ (.A(_03296_),
    .B(_03298_),
    .Y(_03299_));
 sky130_fd_sc_hd__o21ba_1 _23111_ (.A1(_03160_),
    .A2(_03163_),
    .B1_N(_03161_),
    .X(_03300_));
 sky130_fd_sc_hd__o21ba_1 _23112_ (.A1(_03176_),
    .A2(_03180_),
    .B1_N(_03177_),
    .X(_03301_));
 sky130_fd_sc_hd__buf_1 _23113_ (.A(_13739_),
    .X(_03302_));
 sky130_fd_sc_hd__clkbuf_2 _23114_ (.A(_13741_),
    .X(_03303_));
 sky130_fd_sc_hd__a22oi_1 _23115_ (.A1(_14081_),
    .A2(_03302_),
    .B1(_03303_),
    .B2(_13891_),
    .Y(_03304_));
 sky130_fd_sc_hd__and4_1 _23116_ (.A(_14269_),
    .B(_14444_),
    .C(_12772_),
    .D(_13961_),
    .X(_03305_));
 sky130_fd_sc_hd__nor2_1 _23117_ (.A(_03304_),
    .B(_03305_),
    .Y(_03306_));
 sky130_fd_sc_hd__buf_2 _23118_ (.A(_13738_),
    .X(_03307_));
 sky130_fd_sc_hd__buf_2 _23119_ (.A(_13860_),
    .X(_03308_));
 sky130_fd_sc_hd__nand2_1 _23120_ (.A(_03307_),
    .B(_03308_),
    .Y(_03309_));
 sky130_fd_sc_hd__xnor2_1 _23121_ (.A(_03306_),
    .B(_03309_),
    .Y(_03310_));
 sky130_fd_sc_hd__xnor2_1 _23122_ (.A(_03301_),
    .B(_03310_),
    .Y(_03311_));
 sky130_fd_sc_hd__xnor2_1 _23123_ (.A(_03300_),
    .B(_03311_),
    .Y(_03312_));
 sky130_fd_sc_hd__xnor2_1 _23124_ (.A(_03299_),
    .B(_03312_),
    .Y(_03313_));
 sky130_fd_sc_hd__and2b_1 _23125_ (.A_N(_03182_),
    .B(_03184_),
    .X(_03314_));
 sky130_fd_sc_hd__a21oi_1 _23126_ (.A1(_03166_),
    .A2(_03185_),
    .B1(_03314_),
    .Y(_03315_));
 sky130_fd_sc_hd__xor2_1 _23127_ (.A(_03313_),
    .B(_03315_),
    .X(_03316_));
 sky130_fd_sc_hd__xnor2_1 _23128_ (.A(_03280_),
    .B(_03316_),
    .Y(_03317_));
 sky130_fd_sc_hd__and2b_1 _23129_ (.A_N(_03189_),
    .B(_03186_),
    .X(_03318_));
 sky130_fd_sc_hd__a21oi_1 _23130_ (.A1(_03156_),
    .A2(_03190_),
    .B1(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hd__nor2_1 _23131_ (.A(_03317_),
    .B(_03319_),
    .Y(_03320_));
 sky130_fd_sc_hd__and2_1 _23132_ (.A(_03317_),
    .B(_03319_),
    .X(_03321_));
 sky130_fd_sc_hd__or2_1 _23133_ (.A(_03320_),
    .B(_03321_),
    .X(_03322_));
 sky130_fd_sc_hd__xnor2_1 _23134_ (.A(_03259_),
    .B(_03322_),
    .Y(_03323_));
 sky130_fd_sc_hd__nand2_1 _23135_ (.A(_03191_),
    .B(_03193_),
    .Y(_03324_));
 sky130_fd_sc_hd__nor2_1 _23136_ (.A(_03191_),
    .B(_03193_),
    .Y(_03325_));
 sky130_fd_sc_hd__a21oi_1 _23137_ (.A1(_03135_),
    .A2(_03324_),
    .B1(_03325_),
    .Y(_03326_));
 sky130_fd_sc_hd__xnor2_1 _23138_ (.A(_03323_),
    .B(_03326_),
    .Y(_03327_));
 sky130_fd_sc_hd__or2_1 _23139_ (.A(_03237_),
    .B(_03327_),
    .X(_03328_));
 sky130_fd_sc_hd__nand2_1 _23140_ (.A(_03237_),
    .B(_03327_),
    .Y(_03329_));
 sky130_fd_sc_hd__and2_1 _23141_ (.A(_03328_),
    .B(_03329_),
    .X(_03330_));
 sky130_fd_sc_hd__or2_1 _23142_ (.A(_03113_),
    .B(_03198_),
    .X(_03331_));
 sky130_fd_sc_hd__o21ai_2 _23143_ (.A1(_03195_),
    .A2(_03197_),
    .B1(_03331_),
    .Y(_03332_));
 sky130_fd_sc_hd__xor2_1 _23144_ (.A(_03330_),
    .B(_03332_),
    .X(_03333_));
 sky130_fd_sc_hd__xnor2_1 _23145_ (.A(_03222_),
    .B(_03333_),
    .Y(_03334_));
 sky130_fd_sc_hd__and2_1 _23146_ (.A(_03199_),
    .B(_03202_),
    .X(_03335_));
 sky130_fd_sc_hd__or2_1 _23147_ (.A(_03199_),
    .B(_03202_),
    .X(_03336_));
 sky130_fd_sc_hd__o21a_1 _23148_ (.A1(_03098_),
    .A2(_03335_),
    .B1(_03336_),
    .X(_03337_));
 sky130_fd_sc_hd__xnor2_1 _23149_ (.A(_03334_),
    .B(_03337_),
    .Y(_03338_));
 sky130_fd_sc_hd__nand2_1 _23150_ (.A(_03096_),
    .B(_03338_),
    .Y(_03339_));
 sky130_fd_sc_hd__or2_1 _23151_ (.A(_03096_),
    .B(_03338_),
    .X(_03340_));
 sky130_fd_sc_hd__nand2_2 _23152_ (.A(_03339_),
    .B(_03340_),
    .Y(_03341_));
 sky130_fd_sc_hd__nand2_1 _23153_ (.A(_03204_),
    .B(_03207_),
    .Y(_03342_));
 sky130_fd_sc_hd__a21bo_2 _23154_ (.A1(_03093_),
    .A2(_03208_),
    .B1_N(_03342_),
    .X(_03343_));
 sky130_fd_sc_hd__xnor2_4 _23155_ (.A(_03341_),
    .B(_03343_),
    .Y(_03344_));
 sky130_fd_sc_hd__and3b_1 _23156_ (.A_N(_03212_),
    .B(_03087_),
    .C(_03210_),
    .X(_03345_));
 sky130_fd_sc_hd__or3b_2 _23157_ (.A(_02831_),
    .B(_03088_),
    .C_N(_03345_),
    .X(_03346_));
 sky130_fd_sc_hd__nor4_1 _23158_ (.A(_02277_),
    .B(_02420_),
    .C(_02421_),
    .D(_03346_),
    .Y(_03347_));
 sky130_fd_sc_hd__o31ai_4 _23159_ (.A1(_02281_),
    .A2(_02283_),
    .A3(_02284_),
    .B1(net333),
    .Y(_03348_));
 sky130_fd_sc_hd__or3b_1 _23160_ (.A(_02834_),
    .B(_03088_),
    .C_N(_03345_),
    .X(_03349_));
 sky130_fd_sc_hd__or2b_1 _23161_ (.A(_03089_),
    .B_N(_03345_),
    .X(_03350_));
 sky130_fd_sc_hd__o21ai_1 _23162_ (.A1(_03214_),
    .A2(_03212_),
    .B1(_03210_),
    .Y(_03351_));
 sky130_fd_sc_hd__o2111a_2 _23163_ (.A1(_02563_),
    .A2(_03346_),
    .B1(_03349_),
    .C1(_03350_),
    .D1(_03351_),
    .X(_03352_));
 sky130_fd_sc_hd__nand2_2 _23164_ (.A(_03348_),
    .B(_03352_),
    .Y(_03353_));
 sky130_fd_sc_hd__xor2_4 _23165_ (.A(_03344_),
    .B(_03353_),
    .X(_00094_));
 sky130_fd_sc_hd__and3_1 _23166_ (.A(_03339_),
    .B(_03340_),
    .C(_03343_),
    .X(_03354_));
 sky130_fd_sc_hd__a21oi_2 _23167_ (.A1(_03344_),
    .A2(_03353_),
    .B1(_03354_),
    .Y(_03355_));
 sky130_fd_sc_hd__or2b_1 _23168_ (.A(_03337_),
    .B_N(_03334_),
    .X(_03356_));
 sky130_fd_sc_hd__nand2_1 _23169_ (.A(_03226_),
    .B(_03236_),
    .Y(_03357_));
 sky130_fd_sc_hd__a21oi_2 _23170_ (.A1(_03234_),
    .A2(_03357_),
    .B1(_02427_),
    .Y(_03358_));
 sky130_fd_sc_hd__and3_1 _23171_ (.A(_03219_),
    .B(_03234_),
    .C(_03357_),
    .X(_03359_));
 sky130_fd_sc_hd__nor2_1 _23172_ (.A(_03358_),
    .B(_03359_),
    .Y(_03360_));
 sky130_fd_sc_hd__and3_2 _23173_ (.A(_02445_),
    .B(_02853_),
    .C(_03229_),
    .X(_03361_));
 sky130_fd_sc_hd__o21bai_2 _23174_ (.A1(_02433_),
    .A2(_03232_),
    .B1_N(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__and2b_1 _23175_ (.A_N(_03239_),
    .B(_03258_),
    .X(_03363_));
 sky130_fd_sc_hd__nor2_1 _23176_ (.A(_03256_),
    .B(_03363_),
    .Y(_03364_));
 sky130_fd_sc_hd__nor3_2 _23177_ (.A(_02136_),
    .B(_03231_),
    .C(_03361_),
    .Y(_03365_));
 sky130_fd_sc_hd__o21a_1 _23178_ (.A1(_03231_),
    .A2(_03361_),
    .B1(_02136_),
    .X(_03366_));
 sky130_fd_sc_hd__nor2_1 _23179_ (.A(_03365_),
    .B(_03366_),
    .Y(_03367_));
 sky130_fd_sc_hd__buf_2 _23180_ (.A(_03367_),
    .X(_03368_));
 sky130_fd_sc_hd__xnor2_1 _23181_ (.A(_03364_),
    .B(_03368_),
    .Y(_03369_));
 sky130_fd_sc_hd__xnor2_1 _23182_ (.A(_03362_),
    .B(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hd__nor2_1 _23183_ (.A(_03259_),
    .B(_03322_),
    .Y(_03371_));
 sky130_fd_sc_hd__o21ba_1 _23184_ (.A1(_03238_),
    .A2(_03253_),
    .B1_N(_03252_),
    .X(_03372_));
 sky130_vsdinv _23185_ (.A(_03277_),
    .Y(_03373_));
 sky130_fd_sc_hd__or2b_1 _23186_ (.A(_03279_),
    .B_N(_03261_),
    .X(_03374_));
 sky130_fd_sc_hd__o2bb2a_1 _23187_ (.A1_N(_14212_),
    .A2_N(_03245_),
    .B1(_03247_),
    .B2(_03126_),
    .X(_03375_));
 sky130_fd_sc_hd__a31o_1 _23188_ (.A1(_11772_),
    .A2(_14023_),
    .A3(_03266_),
    .B1(_03265_),
    .X(_03376_));
 sky130_fd_sc_hd__o21ai_4 _23189_ (.A1(_14105_),
    .A2(_11782_),
    .B1(_13842_),
    .Y(_03377_));
 sky130_fd_sc_hd__nor2_1 _23190_ (.A(_03245_),
    .B(_03377_),
    .Y(_03378_));
 sky130_fd_sc_hd__xnor2_1 _23191_ (.A(_03126_),
    .B(_03378_),
    .Y(_03379_));
 sky130_fd_sc_hd__clkbuf_2 _23192_ (.A(_03379_),
    .X(_03380_));
 sky130_fd_sc_hd__xor2_1 _23193_ (.A(_03376_),
    .B(_03380_),
    .X(_03381_));
 sky130_fd_sc_hd__and2b_1 _23194_ (.A_N(_03375_),
    .B(_03381_),
    .X(_03382_));
 sky130_fd_sc_hd__and2b_1 _23195_ (.A_N(_03381_),
    .B(_03375_),
    .X(_03383_));
 sky130_fd_sc_hd__or2_1 _23196_ (.A(_03382_),
    .B(_03383_),
    .X(_03384_));
 sky130_fd_sc_hd__and2b_1 _23197_ (.A_N(_03243_),
    .B(_03248_),
    .X(_03385_));
 sky130_fd_sc_hd__and2b_1 _23198_ (.A_N(_03250_),
    .B(_03249_),
    .X(_03386_));
 sky130_fd_sc_hd__nor2_1 _23199_ (.A(_03385_),
    .B(_03386_),
    .Y(_03387_));
 sky130_fd_sc_hd__xor2_1 _23200_ (.A(_03384_),
    .B(_03387_),
    .X(_03388_));
 sky130_fd_sc_hd__xnor2_1 _23201_ (.A(_03240_),
    .B(_03388_),
    .Y(_03389_));
 sky130_fd_sc_hd__a21oi_1 _23202_ (.A1(_03373_),
    .A2(_03374_),
    .B1(_03389_),
    .Y(_03390_));
 sky130_fd_sc_hd__nand3_1 _23203_ (.A(_03373_),
    .B(_03374_),
    .C(_03389_),
    .Y(_03391_));
 sky130_fd_sc_hd__and2b_1 _23204_ (.A_N(_03390_),
    .B(_03391_),
    .X(_03392_));
 sky130_fd_sc_hd__xor2_1 _23205_ (.A(_03372_),
    .B(_03392_),
    .X(_03393_));
 sky130_fd_sc_hd__and2b_2 _23206_ (.A_N(_11819_),
    .B(_01618_),
    .X(_03394_));
 sky130_fd_sc_hd__nand2_2 _23207_ (.A(_11831_),
    .B(_14168_),
    .Y(_03395_));
 sky130_fd_sc_hd__xnor2_4 _23208_ (.A(_03394_),
    .B(_03395_),
    .Y(_03396_));
 sky130_fd_sc_hd__nand2_2 _23209_ (.A(_14457_),
    .B(_14166_),
    .Y(_03397_));
 sky130_fd_sc_hd__xnor2_4 _23210_ (.A(_03396_),
    .B(_03397_),
    .Y(_03398_));
 sky130_fd_sc_hd__and3_1 _23211_ (.A(_12075_),
    .B(_13754_),
    .C(_03281_),
    .X(_03399_));
 sky130_fd_sc_hd__a31o_1 _23212_ (.A1(_14283_),
    .A2(_03286_),
    .A3(_03283_),
    .B1(_03399_),
    .X(_03400_));
 sky130_fd_sc_hd__xor2_2 _23213_ (.A(_03398_),
    .B(_03400_),
    .X(_03401_));
 sky130_fd_sc_hd__clkbuf_2 _23214_ (.A(_13228_),
    .X(_03402_));
 sky130_fd_sc_hd__a22oi_2 _23215_ (.A1(_01564_),
    .A2(_03402_),
    .B1(_03175_),
    .B2(_01558_),
    .Y(_03403_));
 sky130_fd_sc_hd__and4_1 _23216_ (.A(_13667_),
    .B(_13893_),
    .C(_13229_),
    .D(_01613_),
    .X(_03404_));
 sky130_fd_sc_hd__nor2_1 _23217_ (.A(_03403_),
    .B(_03404_),
    .Y(_03405_));
 sky130_fd_sc_hd__nand2_1 _23218_ (.A(_01885_),
    .B(_03179_),
    .Y(_03406_));
 sky130_fd_sc_hd__xnor2_2 _23219_ (.A(_03405_),
    .B(_03406_),
    .Y(_03407_));
 sky130_fd_sc_hd__xnor2_2 _23220_ (.A(_03401_),
    .B(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__and2_1 _23221_ (.A(_03285_),
    .B(_03289_),
    .X(_03409_));
 sky130_fd_sc_hd__a21o_1 _23222_ (.A1(_03290_),
    .A2(_03295_),
    .B1(_03409_),
    .X(_03410_));
 sky130_fd_sc_hd__xnor2_2 _23223_ (.A(_03408_),
    .B(_03410_),
    .Y(_03411_));
 sky130_fd_sc_hd__o21ba_1 _23224_ (.A1(_03304_),
    .A2(_03309_),
    .B1_N(_03305_),
    .X(_03412_));
 sky130_fd_sc_hd__o21ba_1 _23225_ (.A1(_03291_),
    .A2(_03294_),
    .B1_N(_03292_),
    .X(_03413_));
 sky130_fd_sc_hd__a22oi_2 _23226_ (.A1(_14076_),
    .A2(_13739_),
    .B1(_13961_),
    .B2(_13887_),
    .Y(_03414_));
 sky130_fd_sc_hd__and4_1 _23227_ (.A(_14080_),
    .B(_13859_),
    .C(_13743_),
    .D(_13744_),
    .X(_03415_));
 sky130_fd_sc_hd__nor2_1 _23228_ (.A(_03414_),
    .B(_03415_),
    .Y(_03416_));
 sky130_fd_sc_hd__nand2_1 _23229_ (.A(_13738_),
    .B(_14262_),
    .Y(_03417_));
 sky130_fd_sc_hd__xnor2_1 _23230_ (.A(_03416_),
    .B(_03417_),
    .Y(_03418_));
 sky130_fd_sc_hd__xnor2_1 _23231_ (.A(_03413_),
    .B(_03418_),
    .Y(_03419_));
 sky130_fd_sc_hd__xnor2_2 _23232_ (.A(_03412_),
    .B(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__xnor2_2 _23233_ (.A(_03411_),
    .B(_03420_),
    .Y(_03421_));
 sky130_fd_sc_hd__and2b_1 _23234_ (.A_N(_03296_),
    .B(_03298_),
    .X(_03422_));
 sky130_fd_sc_hd__a21oi_2 _23235_ (.A1(_03299_),
    .A2(_03312_),
    .B1(_03422_),
    .Y(_03423_));
 sky130_fd_sc_hd__xor2_2 _23236_ (.A(_03421_),
    .B(_03423_),
    .X(_03424_));
 sky130_fd_sc_hd__or2b_1 _23237_ (.A(_03274_),
    .B_N(_03273_),
    .X(_03425_));
 sky130_fd_sc_hd__a21bo_1 _23238_ (.A1(_03268_),
    .A2(_03275_),
    .B1_N(_03425_),
    .X(_03426_));
 sky130_fd_sc_hd__or2b_1 _23239_ (.A(_03301_),
    .B_N(_03310_),
    .X(_03427_));
 sky130_fd_sc_hd__or2b_1 _23240_ (.A(_03300_),
    .B_N(_03311_),
    .X(_03428_));
 sky130_fd_sc_hd__a22oi_1 _23241_ (.A1(_01757_),
    .A2(_13814_),
    .B1(_13826_),
    .B2(_01582_),
    .Y(_03429_));
 sky130_fd_sc_hd__and4_1 _23242_ (.A(_13936_),
    .B(_01755_),
    .C(_14033_),
    .D(_01846_),
    .X(_03430_));
 sky130_fd_sc_hd__nor2_1 _23243_ (.A(_03429_),
    .B(_03430_),
    .Y(_03431_));
 sky130_fd_sc_hd__nand2_1 _23244_ (.A(_11773_),
    .B(_14212_),
    .Y(_03432_));
 sky130_fd_sc_hd__xnor2_1 _23245_ (.A(_03431_),
    .B(_03432_),
    .Y(_03433_));
 sky130_fd_sc_hd__clkbuf_2 _23246_ (.A(_14310_),
    .X(_03434_));
 sky130_fd_sc_hd__clkbuf_2 _23247_ (.A(_14132_),
    .X(_03435_));
 sky130_fd_sc_hd__a22oi_2 _23248_ (.A1(_03434_),
    .A2(_01538_),
    .B1(_01866_),
    .B2(_03435_),
    .Y(_03436_));
 sky130_fd_sc_hd__and4_1 _23249_ (.A(_12324_),
    .B(_13945_),
    .C(_13868_),
    .D(_01713_),
    .X(_03437_));
 sky130_fd_sc_hd__nor2_1 _23250_ (.A(_03436_),
    .B(_03437_),
    .Y(_03438_));
 sky130_fd_sc_hd__nand2_1 _23251_ (.A(_12228_),
    .B(_01717_),
    .Y(_03439_));
 sky130_fd_sc_hd__xnor2_1 _23252_ (.A(_03438_),
    .B(_03439_),
    .Y(_03440_));
 sky130_fd_sc_hd__o21ba_1 _23253_ (.A1(_03269_),
    .A2(_03272_),
    .B1_N(_03270_),
    .X(_03441_));
 sky130_fd_sc_hd__xnor2_1 _23254_ (.A(_03440_),
    .B(_03441_),
    .Y(_03442_));
 sky130_fd_sc_hd__xnor2_1 _23255_ (.A(_03433_),
    .B(_03442_),
    .Y(_03443_));
 sky130_fd_sc_hd__a21oi_1 _23256_ (.A1(_03427_),
    .A2(_03428_),
    .B1(_03443_),
    .Y(_03444_));
 sky130_fd_sc_hd__and3_1 _23257_ (.A(_03427_),
    .B(_03428_),
    .C(_03443_),
    .X(_03445_));
 sky130_fd_sc_hd__nor2_1 _23258_ (.A(_03444_),
    .B(_03445_),
    .Y(_03446_));
 sky130_fd_sc_hd__xor2_2 _23259_ (.A(_03426_),
    .B(_03446_),
    .X(_03447_));
 sky130_fd_sc_hd__xor2_2 _23260_ (.A(_03424_),
    .B(_03447_),
    .X(_03448_));
 sky130_fd_sc_hd__nor2_1 _23261_ (.A(_03313_),
    .B(_03315_),
    .Y(_03449_));
 sky130_fd_sc_hd__a21o_1 _23262_ (.A1(_03280_),
    .A2(_03316_),
    .B1(_03449_),
    .X(_03450_));
 sky130_fd_sc_hd__xor2_1 _23263_ (.A(_03448_),
    .B(_03450_),
    .X(_03451_));
 sky130_fd_sc_hd__xnor2_1 _23264_ (.A(_03393_),
    .B(_03451_),
    .Y(_03452_));
 sky130_fd_sc_hd__o21a_1 _23265_ (.A1(_03320_),
    .A2(_03371_),
    .B1(_03452_),
    .X(_03453_));
 sky130_fd_sc_hd__nor3_1 _23266_ (.A(_03320_),
    .B(_03371_),
    .C(_03452_),
    .Y(_03454_));
 sky130_fd_sc_hd__nor2_1 _23267_ (.A(_03453_),
    .B(_03454_),
    .Y(_03455_));
 sky130_fd_sc_hd__xnor2_1 _23268_ (.A(_03370_),
    .B(_03455_),
    .Y(_03456_));
 sky130_fd_sc_hd__o21a_1 _23269_ (.A1(_03323_),
    .A2(_03326_),
    .B1(_03328_),
    .X(_03457_));
 sky130_fd_sc_hd__xnor2_1 _23270_ (.A(_03456_),
    .B(_03457_),
    .Y(_03458_));
 sky130_fd_sc_hd__xor2_1 _23271_ (.A(_03360_),
    .B(_03458_),
    .X(_03459_));
 sky130_fd_sc_hd__nor2_1 _23272_ (.A(_03330_),
    .B(_03332_),
    .Y(_03460_));
 sky130_fd_sc_hd__nand2_1 _23273_ (.A(_03330_),
    .B(_03332_),
    .Y(_03461_));
 sky130_fd_sc_hd__o21a_1 _23274_ (.A1(_03222_),
    .A2(_03460_),
    .B1(_03461_),
    .X(_03462_));
 sky130_fd_sc_hd__xnor2_1 _23275_ (.A(_03459_),
    .B(_03462_),
    .Y(_03463_));
 sky130_fd_sc_hd__xnor2_1 _23276_ (.A(_03220_),
    .B(_03463_),
    .Y(_03464_));
 sky130_fd_sc_hd__a21oi_1 _23277_ (.A1(_03356_),
    .A2(_03339_),
    .B1(_03464_),
    .Y(_03465_));
 sky130_fd_sc_hd__nand3_1 _23278_ (.A(_03356_),
    .B(_03339_),
    .C(_03464_),
    .Y(_03466_));
 sky130_fd_sc_hd__and2b_2 _23279_ (.A_N(_03465_),
    .B(_03466_),
    .X(_03467_));
 sky130_fd_sc_hd__xnor2_4 _23280_ (.A(_03355_),
    .B(_03467_),
    .Y(_00095_));
 sky130_fd_sc_hd__nand2_1 _23281_ (.A(_03344_),
    .B(_03467_),
    .Y(_03468_));
 sky130_fd_sc_hd__a21oi_4 _23282_ (.A1(_03348_),
    .A2(_03352_),
    .B1(_03468_),
    .Y(_03469_));
 sky130_fd_sc_hd__o21a_2 _23283_ (.A1(_03354_),
    .A2(_03465_),
    .B1(_03466_),
    .X(_03470_));
 sky130_fd_sc_hd__clkbuf_2 _23284_ (.A(_03365_),
    .X(_03471_));
 sky130_fd_sc_hd__clkbuf_2 _23285_ (.A(_03366_),
    .X(_03472_));
 sky130_fd_sc_hd__or3_1 _23286_ (.A(_03364_),
    .B(_03471_),
    .C(_03472_),
    .X(_03473_));
 sky130_fd_sc_hd__nand2_1 _23287_ (.A(_03362_),
    .B(_03369_),
    .Y(_03474_));
 sky130_fd_sc_hd__a21oi_1 _23288_ (.A1(_03473_),
    .A2(_03474_),
    .B1(_02425_),
    .Y(_03475_));
 sky130_fd_sc_hd__and3_1 _23289_ (.A(_02425_),
    .B(_03473_),
    .C(_03474_),
    .X(_03476_));
 sky130_fd_sc_hd__or2_1 _23290_ (.A(_03475_),
    .B(_03476_),
    .X(_03477_));
 sky130_fd_sc_hd__nor2_4 _23291_ (.A(_03361_),
    .B(_03365_),
    .Y(_03478_));
 sky130_fd_sc_hd__nor3b_1 _23292_ (.A(_03372_),
    .B(_03390_),
    .C_N(_03391_),
    .Y(_03479_));
 sky130_fd_sc_hd__o21ai_1 _23293_ (.A1(_03390_),
    .A2(_03479_),
    .B1(_03368_),
    .Y(_03480_));
 sky130_fd_sc_hd__or3_1 _23294_ (.A(_03367_),
    .B(_03390_),
    .C(_03479_),
    .X(_03481_));
 sky130_fd_sc_hd__and2_1 _23295_ (.A(_03480_),
    .B(_03481_),
    .X(_03482_));
 sky130_fd_sc_hd__xnor2_1 _23296_ (.A(_03478_),
    .B(_03482_),
    .Y(_03483_));
 sky130_fd_sc_hd__and2b_1 _23297_ (.A_N(_11949_),
    .B(_01618_),
    .X(_03484_));
 sky130_fd_sc_hd__nand2_1 _23298_ (.A(_11959_),
    .B(_14168_),
    .Y(_03485_));
 sky130_fd_sc_hd__xnor2_2 _23299_ (.A(_03484_),
    .B(_03485_),
    .Y(_03486_));
 sky130_fd_sc_hd__nand2_1 _23300_ (.A(_13667_),
    .B(_14166_),
    .Y(_03487_));
 sky130_fd_sc_hd__xnor2_2 _23301_ (.A(_03486_),
    .B(_03487_),
    .Y(_03488_));
 sky130_fd_sc_hd__and3_1 _23302_ (.A(_13904_),
    .B(_01625_),
    .C(_03394_),
    .X(_03489_));
 sky130_fd_sc_hd__a31o_1 _23303_ (.A1(_14457_),
    .A2(_03286_),
    .A3(_03396_),
    .B1(_03489_),
    .X(_03490_));
 sky130_fd_sc_hd__xor2_1 _23304_ (.A(_03488_),
    .B(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__a22oi_1 _23305_ (.A1(_13659_),
    .A2(_03402_),
    .B1(_03175_),
    .B2(_13893_),
    .Y(_03492_));
 sky130_fd_sc_hd__and4_1 _23306_ (.A(_13668_),
    .B(_13891_),
    .C(_13229_),
    .D(_01613_),
    .X(_03493_));
 sky130_fd_sc_hd__nor2_1 _23307_ (.A(_03492_),
    .B(_03493_),
    .Y(_03494_));
 sky130_fd_sc_hd__nand2_1 _23308_ (.A(_02036_),
    .B(_03179_),
    .Y(_03495_));
 sky130_fd_sc_hd__xnor2_1 _23309_ (.A(_03494_),
    .B(_03495_),
    .Y(_03496_));
 sky130_fd_sc_hd__xnor2_1 _23310_ (.A(_03491_),
    .B(_03496_),
    .Y(_03497_));
 sky130_fd_sc_hd__and2_1 _23311_ (.A(_03398_),
    .B(_03400_),
    .X(_03498_));
 sky130_fd_sc_hd__a21o_1 _23312_ (.A1(_03401_),
    .A2(_03407_),
    .B1(_03498_),
    .X(_03499_));
 sky130_fd_sc_hd__xnor2_1 _23313_ (.A(_03497_),
    .B(_03499_),
    .Y(_03500_));
 sky130_fd_sc_hd__o21ba_1 _23314_ (.A1(_03414_),
    .A2(_03417_),
    .B1_N(_03415_),
    .X(_03501_));
 sky130_fd_sc_hd__o21ba_1 _23315_ (.A1(_03403_),
    .A2(_03406_),
    .B1_N(_03404_),
    .X(_03502_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _23316_ (.A(_13739_),
    .X(_03503_));
 sky130_fd_sc_hd__a22oi_1 _23317_ (.A1(_03503_),
    .A2(_01540_),
    .B1(_03303_),
    .B2(_01544_),
    .Y(_03504_));
 sky130_fd_sc_hd__and4_1 _23318_ (.A(_14077_),
    .B(_03302_),
    .C(_13861_),
    .D(_03159_),
    .X(_03505_));
 sky130_fd_sc_hd__nor2_1 _23319_ (.A(_03504_),
    .B(_03505_),
    .Y(_03506_));
 sky130_fd_sc_hd__nand2_1 _23320_ (.A(_03307_),
    .B(_13869_),
    .Y(_03507_));
 sky130_fd_sc_hd__xnor2_1 _23321_ (.A(_03506_),
    .B(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__xnor2_1 _23322_ (.A(_03502_),
    .B(_03508_),
    .Y(_03509_));
 sky130_fd_sc_hd__xnor2_1 _23323_ (.A(_03501_),
    .B(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hd__xnor2_1 _23324_ (.A(_03500_),
    .B(_03510_),
    .Y(_03511_));
 sky130_fd_sc_hd__and2b_1 _23325_ (.A_N(_03408_),
    .B(_03410_),
    .X(_03512_));
 sky130_fd_sc_hd__a21oi_1 _23326_ (.A1(_03411_),
    .A2(_03420_),
    .B1(_03512_),
    .Y(_03513_));
 sky130_fd_sc_hd__xor2_1 _23327_ (.A(_03511_),
    .B(_03513_),
    .X(_03514_));
 sky130_fd_sc_hd__and2b_1 _23328_ (.A_N(_03441_),
    .B(_03440_),
    .X(_03515_));
 sky130_fd_sc_hd__a21oi_1 _23329_ (.A1(_03433_),
    .A2(_03442_),
    .B1(_03515_),
    .Y(_03516_));
 sky130_fd_sc_hd__and2b_1 _23330_ (.A_N(_03413_),
    .B(_03418_),
    .X(_03517_));
 sky130_fd_sc_hd__and2b_1 _23331_ (.A_N(_03412_),
    .B(_03419_),
    .X(_03518_));
 sky130_fd_sc_hd__a22oi_2 _23332_ (.A1(_01583_),
    .A2(_13826_),
    .B1(_13831_),
    .B2(_11892_),
    .Y(_03519_));
 sky130_fd_sc_hd__and4_2 _23333_ (.A(_13936_),
    .B(_13937_),
    .C(_14225_),
    .D(_13830_),
    .X(_03520_));
 sky130_fd_sc_hd__nand2_4 _23334_ (.A(_13711_),
    .B(_14570_),
    .Y(_03521_));
 sky130_fd_sc_hd__o21a_1 _23335_ (.A1(_03519_),
    .A2(_03520_),
    .B1(_03521_),
    .X(_03522_));
 sky130_fd_sc_hd__nor3_1 _23336_ (.A(_03519_),
    .B(_03520_),
    .C(_03521_),
    .Y(_03523_));
 sky130_fd_sc_hd__or2_1 _23337_ (.A(_03522_),
    .B(_03523_),
    .X(_03524_));
 sky130_fd_sc_hd__a22oi_2 _23338_ (.A1(_13945_),
    .A2(_13446_),
    .B1(_13836_),
    .B2(_12324_),
    .Y(_03525_));
 sky130_fd_sc_hd__and4_1 _23339_ (.A(_14132_),
    .B(_13721_),
    .C(_13838_),
    .D(_13839_),
    .X(_03526_));
 sky130_fd_sc_hd__nor2_1 _23340_ (.A(_03525_),
    .B(_03526_),
    .Y(_03527_));
 sky130_fd_sc_hd__nand2_1 _23341_ (.A(_12228_),
    .B(_01870_),
    .Y(_03528_));
 sky130_fd_sc_hd__xnor2_1 _23342_ (.A(_03527_),
    .B(_03528_),
    .Y(_03529_));
 sky130_fd_sc_hd__o21ba_1 _23343_ (.A1(_03436_),
    .A2(_03439_),
    .B1_N(_03437_),
    .X(_03530_));
 sky130_fd_sc_hd__xnor2_1 _23344_ (.A(_03529_),
    .B(_03530_),
    .Y(_03531_));
 sky130_fd_sc_hd__xnor2_1 _23345_ (.A(_03524_),
    .B(_03531_),
    .Y(_03532_));
 sky130_fd_sc_hd__o21a_1 _23346_ (.A1(_03517_),
    .A2(_03518_),
    .B1(_03532_),
    .X(_03533_));
 sky130_fd_sc_hd__or3_1 _23347_ (.A(_03517_),
    .B(_03518_),
    .C(_03532_),
    .X(_03534_));
 sky130_fd_sc_hd__and2b_1 _23348_ (.A_N(_03533_),
    .B(_03534_),
    .X(_03535_));
 sky130_fd_sc_hd__xnor2_1 _23349_ (.A(_03516_),
    .B(_03535_),
    .Y(_03536_));
 sky130_fd_sc_hd__xnor2_1 _23350_ (.A(_03514_),
    .B(_03536_),
    .Y(_03537_));
 sky130_fd_sc_hd__nor2_1 _23351_ (.A(_03421_),
    .B(_03423_),
    .Y(_03538_));
 sky130_fd_sc_hd__a21oi_1 _23352_ (.A1(_03424_),
    .A2(_03447_),
    .B1(_03538_),
    .Y(_03539_));
 sky130_fd_sc_hd__nor2_1 _23353_ (.A(_03537_),
    .B(_03539_),
    .Y(_03540_));
 sky130_fd_sc_hd__and2_1 _23354_ (.A(_03537_),
    .B(_03539_),
    .X(_03541_));
 sky130_fd_sc_hd__or2_1 _23355_ (.A(_03540_),
    .B(_03541_),
    .X(_03542_));
 sky130_fd_sc_hd__nor2_1 _23356_ (.A(_03384_),
    .B(_03387_),
    .Y(_03543_));
 sky130_fd_sc_hd__and2_1 _23357_ (.A(_03240_),
    .B(_03388_),
    .X(_03544_));
 sky130_fd_sc_hd__a21oi_1 _23358_ (.A1(_03426_),
    .A2(_03446_),
    .B1(_03444_),
    .Y(_03545_));
 sky130_fd_sc_hd__and2_1 _23359_ (.A(_03376_),
    .B(_03380_),
    .X(_03546_));
 sky130_fd_sc_hd__clkbuf_2 _23360_ (.A(_13827_),
    .X(_03547_));
 sky130_fd_sc_hd__a31o_1 _23361_ (.A1(_11772_),
    .A2(_03547_),
    .A3(_03431_),
    .B1(_03430_),
    .X(_03548_));
 sky130_fd_sc_hd__xor2_1 _23362_ (.A(_03379_),
    .B(_03548_),
    .X(_03549_));
 sky130_fd_sc_hd__a21oi_2 _23363_ (.A1(_03244_),
    .A2(_03378_),
    .B1(_03245_),
    .Y(_03550_));
 sky130_fd_sc_hd__xnor2_1 _23364_ (.A(_03549_),
    .B(_03550_),
    .Y(_03551_));
 sky130_fd_sc_hd__o21a_1 _23365_ (.A1(_03546_),
    .A2(_03382_),
    .B1(_03551_),
    .X(_03552_));
 sky130_fd_sc_hd__nor3_1 _23366_ (.A(_03546_),
    .B(_03382_),
    .C(_03551_),
    .Y(_03553_));
 sky130_fd_sc_hd__nor2_1 _23367_ (.A(_03552_),
    .B(_03553_),
    .Y(_03554_));
 sky130_fd_sc_hd__xnor2_1 _23368_ (.A(_03118_),
    .B(_03554_),
    .Y(_03555_));
 sky130_fd_sc_hd__xnor2_1 _23369_ (.A(_03545_),
    .B(_03555_),
    .Y(_03556_));
 sky130_fd_sc_hd__o21a_1 _23370_ (.A1(_03543_),
    .A2(_03544_),
    .B1(_03556_),
    .X(_03557_));
 sky130_fd_sc_hd__nor3_1 _23371_ (.A(_03543_),
    .B(_03544_),
    .C(_03556_),
    .Y(_03558_));
 sky130_fd_sc_hd__or2_1 _23372_ (.A(_03557_),
    .B(_03558_),
    .X(_03559_));
 sky130_fd_sc_hd__xor2_1 _23373_ (.A(_03542_),
    .B(_03559_),
    .X(_03560_));
 sky130_fd_sc_hd__nor2_1 _23374_ (.A(_03448_),
    .B(_03450_),
    .Y(_03561_));
 sky130_fd_sc_hd__nand2_1 _23375_ (.A(_03448_),
    .B(_03450_),
    .Y(_03562_));
 sky130_fd_sc_hd__o21a_1 _23376_ (.A1(_03393_),
    .A2(_03561_),
    .B1(_03562_),
    .X(_03563_));
 sky130_fd_sc_hd__xnor2_1 _23377_ (.A(_03560_),
    .B(_03563_),
    .Y(_03564_));
 sky130_fd_sc_hd__xor2_1 _23378_ (.A(_03483_),
    .B(_03564_),
    .X(_03565_));
 sky130_fd_sc_hd__o21ba_1 _23379_ (.A1(_03370_),
    .A2(_03454_),
    .B1_N(_03453_),
    .X(_03566_));
 sky130_fd_sc_hd__xor2_1 _23380_ (.A(_03565_),
    .B(_03566_),
    .X(_03567_));
 sky130_fd_sc_hd__nor2_1 _23381_ (.A(_03477_),
    .B(_03567_),
    .Y(_03568_));
 sky130_fd_sc_hd__and2_1 _23382_ (.A(_03477_),
    .B(_03567_),
    .X(_03569_));
 sky130_fd_sc_hd__or2_1 _23383_ (.A(_03568_),
    .B(_03569_),
    .X(_03570_));
 sky130_fd_sc_hd__or2b_1 _23384_ (.A(_03457_),
    .B_N(_03456_),
    .X(_03571_));
 sky130_fd_sc_hd__a21bo_1 _23385_ (.A1(_03360_),
    .A2(_03458_),
    .B1_N(_03571_),
    .X(_03572_));
 sky130_fd_sc_hd__xnor2_1 _23386_ (.A(_03570_),
    .B(_03572_),
    .Y(_03573_));
 sky130_fd_sc_hd__xnor2_1 _23387_ (.A(_03358_),
    .B(_03573_),
    .Y(_03574_));
 sky130_fd_sc_hd__or2b_1 _23388_ (.A(_03462_),
    .B_N(_03459_),
    .X(_03575_));
 sky130_fd_sc_hd__a21bo_1 _23389_ (.A1(_03220_),
    .A2(_03463_),
    .B1_N(_03575_),
    .X(_03576_));
 sky130_fd_sc_hd__xnor2_1 _23390_ (.A(_03574_),
    .B(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hd__o21a_1 _23391_ (.A1(_03469_),
    .A2(_03470_),
    .B1(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__nor3_1 _23392_ (.A(_03577_),
    .B(_03469_),
    .C(_03470_),
    .Y(_03579_));
 sky130_fd_sc_hd__nor2_2 _23393_ (.A(_03578_),
    .B(_03579_),
    .Y(_00096_));
 sky130_fd_sc_hd__or2b_1 _23394_ (.A(_03570_),
    .B_N(_03572_),
    .X(_03580_));
 sky130_fd_sc_hd__nand2_1 _23395_ (.A(_03358_),
    .B(_03573_),
    .Y(_03581_));
 sky130_fd_sc_hd__and2b_1 _23396_ (.A_N(_03566_),
    .B(_03565_),
    .X(_03582_));
 sky130_fd_sc_hd__or2_2 _23397_ (.A(_03361_),
    .B(_03365_),
    .X(_03583_));
 sky130_fd_sc_hd__nand2_1 _23398_ (.A(_03583_),
    .B(_03482_),
    .Y(_03584_));
 sky130_fd_sc_hd__a21oi_1 _23399_ (.A1(_03480_),
    .A2(_03584_),
    .B1(_02425_),
    .Y(_03585_));
 sky130_fd_sc_hd__and3_1 _23400_ (.A(_02425_),
    .B(_03480_),
    .C(_03584_),
    .X(_03586_));
 sky130_fd_sc_hd__or2_1 _23401_ (.A(_03585_),
    .B(_03586_),
    .X(_03587_));
 sky130_fd_sc_hd__and2b_1 _23402_ (.A_N(_12070_),
    .B(_13803_),
    .X(_03588_));
 sky130_fd_sc_hd__nand2_1 _23403_ (.A(_13666_),
    .B(_13757_),
    .Y(_03589_));
 sky130_fd_sc_hd__xnor2_2 _23404_ (.A(_03588_),
    .B(_03589_),
    .Y(_03590_));
 sky130_fd_sc_hd__nand2_1 _23405_ (.A(_13893_),
    .B(_01624_),
    .Y(_03591_));
 sky130_fd_sc_hd__xnor2_2 _23406_ (.A(_03590_),
    .B(_03591_),
    .Y(_03592_));
 sky130_fd_sc_hd__and3_1 _23407_ (.A(_12278_),
    .B(_13754_),
    .C(_03484_),
    .X(_03593_));
 sky130_fd_sc_hd__a31o_1 _23408_ (.A1(_01558_),
    .A2(_03286_),
    .A3(_03486_),
    .B1(_03593_),
    .X(_03594_));
 sky130_fd_sc_hd__xor2_2 _23409_ (.A(_03592_),
    .B(_03594_),
    .X(_03595_));
 sky130_fd_sc_hd__clkbuf_2 _23410_ (.A(_13224_),
    .X(_03596_));
 sky130_fd_sc_hd__clkbuf_2 _23411_ (.A(_14510_),
    .X(_03597_));
 sky130_fd_sc_hd__a22oi_1 _23412_ (.A1(_13888_),
    .A2(_03596_),
    .B1(_03597_),
    .B2(_13659_),
    .Y(_03598_));
 sky130_fd_sc_hd__and4_1 _23413_ (.A(_13659_),
    .B(_14081_),
    .C(_03402_),
    .D(_01613_),
    .X(_03599_));
 sky130_fd_sc_hd__nor2_1 _23414_ (.A(_03598_),
    .B(_03599_),
    .Y(_03600_));
 sky130_fd_sc_hd__nand2_1 _23415_ (.A(_03308_),
    .B(_03179_),
    .Y(_03601_));
 sky130_fd_sc_hd__xnor2_2 _23416_ (.A(_03600_),
    .B(_03601_),
    .Y(_03602_));
 sky130_fd_sc_hd__xnor2_2 _23417_ (.A(_03595_),
    .B(_03602_),
    .Y(_03603_));
 sky130_fd_sc_hd__and2_1 _23418_ (.A(_03488_),
    .B(_03490_),
    .X(_03604_));
 sky130_fd_sc_hd__a21o_1 _23419_ (.A1(_03491_),
    .A2(_03496_),
    .B1(_03604_),
    .X(_03605_));
 sky130_fd_sc_hd__xnor2_1 _23420_ (.A(_03603_),
    .B(_03605_),
    .Y(_03606_));
 sky130_fd_sc_hd__o21ba_1 _23421_ (.A1(_03504_),
    .A2(_03507_),
    .B1_N(_03505_),
    .X(_03607_));
 sky130_fd_sc_hd__o21ba_1 _23422_ (.A1(_03492_),
    .A2(_03495_),
    .B1_N(_03493_),
    .X(_03608_));
 sky130_fd_sc_hd__clkbuf_4 _23423_ (.A(_13961_),
    .X(_03609_));
 sky130_fd_sc_hd__a22oi_1 _23424_ (.A1(_01540_),
    .A2(_03609_),
    .B1(_13869_),
    .B2(_03503_),
    .Y(_03610_));
 sky130_fd_sc_hd__and4_1 _23425_ (.A(_03302_),
    .B(_14262_),
    .C(_03159_),
    .D(_01538_),
    .X(_03611_));
 sky130_fd_sc_hd__nor2_1 _23426_ (.A(_03610_),
    .B(_03611_),
    .Y(_03612_));
 sky130_fd_sc_hd__nand2_1 _23427_ (.A(_12587_),
    .B(_02610_),
    .Y(_03613_));
 sky130_fd_sc_hd__xnor2_1 _23428_ (.A(_03612_),
    .B(_03613_),
    .Y(_03614_));
 sky130_fd_sc_hd__xnor2_1 _23429_ (.A(_03608_),
    .B(_03614_),
    .Y(_03615_));
 sky130_fd_sc_hd__xnor2_1 _23430_ (.A(_03607_),
    .B(_03615_),
    .Y(_03616_));
 sky130_fd_sc_hd__xnor2_1 _23431_ (.A(_03606_),
    .B(_03616_),
    .Y(_03617_));
 sky130_fd_sc_hd__and2b_1 _23432_ (.A_N(_03497_),
    .B(_03499_),
    .X(_03618_));
 sky130_fd_sc_hd__a21oi_1 _23433_ (.A1(_03500_),
    .A2(_03510_),
    .B1(_03618_),
    .Y(_03619_));
 sky130_fd_sc_hd__nor2_1 _23434_ (.A(_03617_),
    .B(_03619_),
    .Y(_03620_));
 sky130_fd_sc_hd__nand2_1 _23435_ (.A(_03617_),
    .B(_03619_),
    .Y(_03621_));
 sky130_fd_sc_hd__or2b_1 _23436_ (.A(_03620_),
    .B_N(_03621_),
    .X(_03622_));
 sky130_fd_sc_hd__or2b_1 _23437_ (.A(_03530_),
    .B_N(_03529_),
    .X(_03623_));
 sky130_fd_sc_hd__or2b_1 _23438_ (.A(_03524_),
    .B_N(_03531_),
    .X(_03624_));
 sky130_fd_sc_hd__nand2_1 _23439_ (.A(_03623_),
    .B(_03624_),
    .Y(_03625_));
 sky130_fd_sc_hd__or2b_1 _23440_ (.A(_03502_),
    .B_N(_03508_),
    .X(_03626_));
 sky130_fd_sc_hd__or2b_1 _23441_ (.A(_03501_),
    .B_N(_03509_),
    .X(_03627_));
 sky130_fd_sc_hd__clkbuf_2 _23442_ (.A(_03547_),
    .X(_03628_));
 sky130_fd_sc_hd__and3_1 _23443_ (.A(_11892_),
    .B(_01583_),
    .C(_14570_),
    .X(_03629_));
 sky130_fd_sc_hd__a22o_1 _23444_ (.A1(_01583_),
    .A2(_03547_),
    .B1(_14038_),
    .B2(_11892_),
    .X(_03630_));
 sky130_fd_sc_hd__a21bo_1 _23445_ (.A1(_03628_),
    .A2(_03629_),
    .B1_N(_03630_),
    .X(_03631_));
 sky130_fd_sc_hd__xor2_1 _23446_ (.A(_03521_),
    .B(_03631_),
    .X(_03632_));
 sky130_fd_sc_hd__clkbuf_4 _23447_ (.A(_13945_),
    .X(_03633_));
 sky130_fd_sc_hd__a22oi_1 _23448_ (.A1(_03633_),
    .A2(_01844_),
    .B1(_13825_),
    .B2(_12325_),
    .Y(_03634_));
 sky130_fd_sc_hd__and4_1 _23449_ (.A(_03435_),
    .B(_03434_),
    .C(_01844_),
    .D(_13825_),
    .X(_03635_));
 sky130_fd_sc_hd__nor2_1 _23450_ (.A(_03634_),
    .B(_03635_),
    .Y(_03636_));
 sky130_fd_sc_hd__nand2_1 _23451_ (.A(_12229_),
    .B(_14023_),
    .Y(_03637_));
 sky130_fd_sc_hd__xnor2_1 _23452_ (.A(_03636_),
    .B(_03637_),
    .Y(_03638_));
 sky130_fd_sc_hd__o21ba_1 _23453_ (.A1(_03525_),
    .A2(_03528_),
    .B1_N(_03526_),
    .X(_03639_));
 sky130_fd_sc_hd__xnor2_1 _23454_ (.A(_03638_),
    .B(_03639_),
    .Y(_03640_));
 sky130_fd_sc_hd__xnor2_1 _23455_ (.A(_03632_),
    .B(_03640_),
    .Y(_03641_));
 sky130_fd_sc_hd__a21o_1 _23456_ (.A1(_03626_),
    .A2(_03627_),
    .B1(_03641_),
    .X(_03642_));
 sky130_fd_sc_hd__nand3_1 _23457_ (.A(_03626_),
    .B(_03627_),
    .C(_03641_),
    .Y(_03643_));
 sky130_fd_sc_hd__nand2_1 _23458_ (.A(_03642_),
    .B(_03643_),
    .Y(_03644_));
 sky130_fd_sc_hd__xnor2_1 _23459_ (.A(_03625_),
    .B(_03644_),
    .Y(_03645_));
 sky130_fd_sc_hd__xnor2_1 _23460_ (.A(_03622_),
    .B(_03645_),
    .Y(_03646_));
 sky130_fd_sc_hd__nor2_1 _23461_ (.A(_03511_),
    .B(_03513_),
    .Y(_03647_));
 sky130_fd_sc_hd__a21o_1 _23462_ (.A1(_03514_),
    .A2(_03536_),
    .B1(_03647_),
    .X(_03648_));
 sky130_fd_sc_hd__xnor2_1 _23463_ (.A(_03646_),
    .B(_03648_),
    .Y(_03649_));
 sky130_fd_sc_hd__a21oi_1 _23464_ (.A1(_03240_),
    .A2(_03554_),
    .B1(_03552_),
    .Y(_03650_));
 sky130_fd_sc_hd__and2b_1 _23465_ (.A_N(_03516_),
    .B(_03535_),
    .X(_03651_));
 sky130_fd_sc_hd__o21a_1 _23466_ (.A1(_03520_),
    .A2(_03523_),
    .B1(_03380_),
    .X(_03652_));
 sky130_fd_sc_hd__nor3_1 _23467_ (.A(_03380_),
    .B(_03520_),
    .C(_03523_),
    .Y(_03653_));
 sky130_fd_sc_hd__nor2_1 _23468_ (.A(_03652_),
    .B(_03653_),
    .Y(_03654_));
 sky130_fd_sc_hd__xnor2_1 _23469_ (.A(_03550_),
    .B(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__nor2_1 _23470_ (.A(_03380_),
    .B(_03548_),
    .Y(_03656_));
 sky130_fd_sc_hd__nand2_1 _23471_ (.A(_03380_),
    .B(_03548_),
    .Y(_03657_));
 sky130_fd_sc_hd__o21a_1 _23472_ (.A1(_03656_),
    .A2(_03550_),
    .B1(_03657_),
    .X(_03658_));
 sky130_fd_sc_hd__xnor2_1 _23473_ (.A(_03655_),
    .B(_03658_),
    .Y(_03659_));
 sky130_fd_sc_hd__xnor2_1 _23474_ (.A(_03118_),
    .B(_03659_),
    .Y(_03660_));
 sky130_fd_sc_hd__o21a_1 _23475_ (.A1(_03533_),
    .A2(_03651_),
    .B1(_03660_),
    .X(_03661_));
 sky130_fd_sc_hd__nor3_1 _23476_ (.A(_03533_),
    .B(_03651_),
    .C(_03660_),
    .Y(_03662_));
 sky130_fd_sc_hd__nor2_1 _23477_ (.A(_03661_),
    .B(_03662_),
    .Y(_03663_));
 sky130_fd_sc_hd__xnor2_1 _23478_ (.A(_03650_),
    .B(_03663_),
    .Y(_03664_));
 sky130_fd_sc_hd__xnor2_1 _23479_ (.A(_03649_),
    .B(_03664_),
    .Y(_03665_));
 sky130_fd_sc_hd__o21ba_1 _23480_ (.A1(_03542_),
    .A2(_03559_),
    .B1_N(_03540_),
    .X(_03666_));
 sky130_fd_sc_hd__xnor2_1 _23481_ (.A(_03665_),
    .B(_03666_),
    .Y(_03667_));
 sky130_fd_sc_hd__and2b_1 _23482_ (.A_N(_03545_),
    .B(_03555_),
    .X(_03668_));
 sky130_fd_sc_hd__o21ai_1 _23483_ (.A1(_03668_),
    .A2(_03557_),
    .B1(_03368_),
    .Y(_03669_));
 sky130_fd_sc_hd__or3_1 _23484_ (.A(_03367_),
    .B(_03668_),
    .C(_03557_),
    .X(_03670_));
 sky130_fd_sc_hd__and2_1 _23485_ (.A(_03669_),
    .B(_03670_),
    .X(_03671_));
 sky130_fd_sc_hd__xnor2_1 _23486_ (.A(_03478_),
    .B(_03671_),
    .Y(_03672_));
 sky130_fd_sc_hd__xnor2_1 _23487_ (.A(_03667_),
    .B(_03672_),
    .Y(_03673_));
 sky130_fd_sc_hd__and2b_1 _23488_ (.A_N(_03563_),
    .B(_03560_),
    .X(_03674_));
 sky130_fd_sc_hd__a21oi_1 _23489_ (.A1(_03483_),
    .A2(_03564_),
    .B1(_03674_),
    .Y(_03675_));
 sky130_fd_sc_hd__nor2_1 _23490_ (.A(_03673_),
    .B(_03675_),
    .Y(_03676_));
 sky130_fd_sc_hd__and2_1 _23491_ (.A(_03673_),
    .B(_03675_),
    .X(_03677_));
 sky130_fd_sc_hd__nor2_1 _23492_ (.A(_03676_),
    .B(_03677_),
    .Y(_03678_));
 sky130_fd_sc_hd__xnor2_1 _23493_ (.A(_03587_),
    .B(_03678_),
    .Y(_03679_));
 sky130_fd_sc_hd__o21ai_1 _23494_ (.A1(_03582_),
    .A2(_03568_),
    .B1(_03679_),
    .Y(_03680_));
 sky130_fd_sc_hd__or3_1 _23495_ (.A(_03582_),
    .B(_03568_),
    .C(_03679_),
    .X(_03681_));
 sky130_fd_sc_hd__and2_1 _23496_ (.A(_03680_),
    .B(_03681_),
    .X(_03682_));
 sky130_fd_sc_hd__xnor2_1 _23497_ (.A(_03475_),
    .B(_03682_),
    .Y(_03683_));
 sky130_fd_sc_hd__and3_1 _23498_ (.A(_03580_),
    .B(_03581_),
    .C(_03683_),
    .X(_03684_));
 sky130_fd_sc_hd__a21oi_1 _23499_ (.A1(_03580_),
    .A2(_03581_),
    .B1(_03683_),
    .Y(_03685_));
 sky130_fd_sc_hd__nor2_2 _23500_ (.A(_03684_),
    .B(_03685_),
    .Y(_03686_));
 sky130_fd_sc_hd__and2b_1 _23501_ (.A_N(_03574_),
    .B(_03576_),
    .X(_03687_));
 sky130_fd_sc_hd__nor2_2 _23502_ (.A(_03687_),
    .B(_03578_),
    .Y(_03688_));
 sky130_fd_sc_hd__xnor2_4 _23503_ (.A(_03686_),
    .B(_03688_),
    .Y(_00097_));
 sky130_fd_sc_hd__nand2_1 _23504_ (.A(_03475_),
    .B(_03682_),
    .Y(_03689_));
 sky130_fd_sc_hd__and2b_1 _23505_ (.A_N(_13663_),
    .B(_13804_),
    .X(_03690_));
 sky130_fd_sc_hd__nand2_1 _23506_ (.A(_13893_),
    .B(_13754_),
    .Y(_03691_));
 sky130_fd_sc_hd__xnor2_2 _23507_ (.A(_03690_),
    .B(_03691_),
    .Y(_03692_));
 sky130_fd_sc_hd__nand2_1 _23508_ (.A(_01885_),
    .B(_03286_),
    .Y(_03693_));
 sky130_fd_sc_hd__xnor2_2 _23509_ (.A(_03692_),
    .B(_03693_),
    .Y(_03694_));
 sky130_fd_sc_hd__buf_2 _23510_ (.A(_01624_),
    .X(_03695_));
 sky130_fd_sc_hd__and3_1 _23511_ (.A(_01558_),
    .B(_03287_),
    .C(_03588_),
    .X(_03696_));
 sky130_fd_sc_hd__a31o_1 _23512_ (.A1(_01564_),
    .A2(_03695_),
    .A3(_03590_),
    .B1(_03696_),
    .X(_03697_));
 sky130_fd_sc_hd__xor2_2 _23513_ (.A(_03694_),
    .B(_03697_),
    .X(_03698_));
 sky130_fd_sc_hd__a22oi_1 _23514_ (.A1(_03308_),
    .A2(_03596_),
    .B1(_03597_),
    .B2(_02036_),
    .Y(_03699_));
 sky130_fd_sc_hd__and4_1 _23515_ (.A(_13888_),
    .B(_01544_),
    .C(_03596_),
    .D(_03597_),
    .X(_03700_));
 sky130_fd_sc_hd__nor2_1 _23516_ (.A(_03699_),
    .B(_03700_),
    .Y(_03701_));
 sky130_fd_sc_hd__nand2_1 _23517_ (.A(_02331_),
    .B(_03179_),
    .Y(_03702_));
 sky130_fd_sc_hd__xnor2_2 _23518_ (.A(_03701_),
    .B(_03702_),
    .Y(_03703_));
 sky130_fd_sc_hd__xnor2_2 _23519_ (.A(_03698_),
    .B(_03703_),
    .Y(_03704_));
 sky130_fd_sc_hd__and2_1 _23520_ (.A(_03592_),
    .B(_03594_),
    .X(_03705_));
 sky130_fd_sc_hd__a21o_1 _23521_ (.A1(_03595_),
    .A2(_03602_),
    .B1(_03705_),
    .X(_03706_));
 sky130_fd_sc_hd__xnor2_1 _23522_ (.A(_03704_),
    .B(_03706_),
    .Y(_03707_));
 sky130_fd_sc_hd__o21ba_1 _23523_ (.A1(_03610_),
    .A2(_03613_),
    .B1_N(_03611_),
    .X(_03708_));
 sky130_fd_sc_hd__o21ba_1 _23524_ (.A1(_03598_),
    .A2(_03601_),
    .B1_N(_03599_),
    .X(_03709_));
 sky130_fd_sc_hd__a22oi_1 _23525_ (.A1(_03303_),
    .A2(_14438_),
    .B1(_14059_),
    .B2(_03503_),
    .Y(_03710_));
 sky130_fd_sc_hd__and4_1 _23526_ (.A(_03302_),
    .B(_03159_),
    .C(_13286_),
    .D(_01866_),
    .X(_03711_));
 sky130_fd_sc_hd__nor2_1 _23527_ (.A(_03710_),
    .B(_03711_),
    .Y(_03712_));
 sky130_fd_sc_hd__nand2_1 _23528_ (.A(_03307_),
    .B(_01718_),
    .Y(_03713_));
 sky130_fd_sc_hd__xnor2_1 _23529_ (.A(_03712_),
    .B(_03713_),
    .Y(_03714_));
 sky130_fd_sc_hd__xnor2_1 _23530_ (.A(_03709_),
    .B(_03714_),
    .Y(_03715_));
 sky130_fd_sc_hd__xnor2_1 _23531_ (.A(_03708_),
    .B(_03715_),
    .Y(_03716_));
 sky130_fd_sc_hd__xnor2_1 _23532_ (.A(_03707_),
    .B(_03716_),
    .Y(_03717_));
 sky130_fd_sc_hd__and2b_1 _23533_ (.A_N(_03603_),
    .B(_03605_),
    .X(_03718_));
 sky130_fd_sc_hd__a21oi_1 _23534_ (.A1(_03606_),
    .A2(_03616_),
    .B1(_03718_),
    .Y(_03719_));
 sky130_fd_sc_hd__xor2_1 _23535_ (.A(_03717_),
    .B(_03719_),
    .X(_03720_));
 sky130_fd_sc_hd__and2b_1 _23536_ (.A_N(_03639_),
    .B(_03638_),
    .X(_03721_));
 sky130_fd_sc_hd__a21oi_1 _23537_ (.A1(_03632_),
    .A2(_03640_),
    .B1(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__or2b_1 _23538_ (.A(_03608_),
    .B_N(_03614_),
    .X(_03723_));
 sky130_fd_sc_hd__or2b_1 _23539_ (.A(_03607_),
    .B_N(_03615_),
    .X(_03724_));
 sky130_fd_sc_hd__or2_1 _23540_ (.A(_01582_),
    .B(_01757_),
    .X(_03725_));
 sky130_fd_sc_hd__and3b_1 _23541_ (.A_N(_03629_),
    .B(_03725_),
    .C(_14562_),
    .X(_03726_));
 sky130_fd_sc_hd__xnor2_4 _23542_ (.A(_03521_),
    .B(_03726_),
    .Y(_03727_));
 sky130_fd_sc_hd__a22oi_2 _23543_ (.A1(_03434_),
    .A2(_13825_),
    .B1(_13817_),
    .B2(_03435_),
    .Y(_03728_));
 sky130_fd_sc_hd__and4_1 _23544_ (.A(_03435_),
    .B(_03434_),
    .C(_01870_),
    .D(_13826_),
    .X(_03729_));
 sky130_fd_sc_hd__nor2_1 _23545_ (.A(_03728_),
    .B(_03729_),
    .Y(_03730_));
 sky130_fd_sc_hd__nand2_1 _23546_ (.A(_12229_),
    .B(_03547_),
    .Y(_03731_));
 sky130_fd_sc_hd__xnor2_1 _23547_ (.A(_03730_),
    .B(_03731_),
    .Y(_03732_));
 sky130_fd_sc_hd__o21ba_1 _23548_ (.A1(_03634_),
    .A2(_03637_),
    .B1_N(_03635_),
    .X(_03733_));
 sky130_fd_sc_hd__xnor2_1 _23549_ (.A(_03732_),
    .B(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__xnor2_1 _23550_ (.A(_03727_),
    .B(_03734_),
    .Y(_03735_));
 sky130_fd_sc_hd__a21o_1 _23551_ (.A1(_03723_),
    .A2(_03724_),
    .B1(_03735_),
    .X(_03736_));
 sky130_fd_sc_hd__nand3_1 _23552_ (.A(_03723_),
    .B(_03724_),
    .C(_03735_),
    .Y(_03737_));
 sky130_fd_sc_hd__and2_1 _23553_ (.A(_03736_),
    .B(_03737_),
    .X(_03738_));
 sky130_fd_sc_hd__xnor2_1 _23554_ (.A(_03722_),
    .B(_03738_),
    .Y(_03739_));
 sky130_fd_sc_hd__xnor2_1 _23555_ (.A(_03720_),
    .B(_03739_),
    .Y(_03740_));
 sky130_fd_sc_hd__a21oi_1 _23556_ (.A1(_03621_),
    .A2(_03645_),
    .B1(_03620_),
    .Y(_03741_));
 sky130_fd_sc_hd__nor2_1 _23557_ (.A(_03740_),
    .B(_03741_),
    .Y(_03742_));
 sky130_fd_sc_hd__and2_1 _23558_ (.A(_03740_),
    .B(_03741_),
    .X(_03743_));
 sky130_fd_sc_hd__nor2_1 _23559_ (.A(_03742_),
    .B(_03743_),
    .Y(_03744_));
 sky130_fd_sc_hd__and2b_1 _23560_ (.A_N(_03658_),
    .B(_03655_),
    .X(_03745_));
 sky130_fd_sc_hd__a21oi_1 _23561_ (.A1(_03240_),
    .A2(_03659_),
    .B1(_03745_),
    .Y(_03746_));
 sky130_fd_sc_hd__a21bo_1 _23562_ (.A1(_03625_),
    .A2(_03643_),
    .B1_N(_03642_),
    .X(_03747_));
 sky130_fd_sc_hd__o21bai_1 _23563_ (.A1(_03550_),
    .A2(_03653_),
    .B1_N(_03652_),
    .Y(_03748_));
 sky130_fd_sc_hd__o2bb2a_1 _23564_ (.A1_N(_14213_),
    .A2_N(_03629_),
    .B1(_03631_),
    .B2(_03521_),
    .X(_03749_));
 sky130_fd_sc_hd__and2_1 _23565_ (.A(_11447_),
    .B(_03245_),
    .X(_03750_));
 sky130_fd_sc_hd__a21o_1 _23566_ (.A1(_03126_),
    .A2(_03377_),
    .B1(_03750_),
    .X(_03751_));
 sky130_fd_sc_hd__xor2_1 _23567_ (.A(_03749_),
    .B(_03751_),
    .X(_03752_));
 sky130_fd_sc_hd__xnor2_1 _23568_ (.A(_03748_),
    .B(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__xnor2_1 _23569_ (.A(_03238_),
    .B(_03753_),
    .Y(_03754_));
 sky130_fd_sc_hd__xnor2_1 _23570_ (.A(_03747_),
    .B(_03754_),
    .Y(_03755_));
 sky130_fd_sc_hd__xnor2_1 _23571_ (.A(_03746_),
    .B(_03755_),
    .Y(_03756_));
 sky130_fd_sc_hd__xnor2_1 _23572_ (.A(_03744_),
    .B(_03756_),
    .Y(_03757_));
 sky130_fd_sc_hd__or2_1 _23573_ (.A(_03646_),
    .B(_03648_),
    .X(_03758_));
 sky130_fd_sc_hd__and2_1 _23574_ (.A(_03646_),
    .B(_03648_),
    .X(_03759_));
 sky130_fd_sc_hd__a21oi_1 _23575_ (.A1(_03758_),
    .A2(_03664_),
    .B1(_03759_),
    .Y(_03760_));
 sky130_fd_sc_hd__nor2_1 _23576_ (.A(_03757_),
    .B(_03760_),
    .Y(_03761_));
 sky130_fd_sc_hd__and2_1 _23577_ (.A(_03757_),
    .B(_03760_),
    .X(_03762_));
 sky130_fd_sc_hd__nor2_1 _23578_ (.A(_03761_),
    .B(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__buf_2 _23579_ (.A(_03368_),
    .X(_03764_));
 sky130_fd_sc_hd__and2b_1 _23580_ (.A_N(_03650_),
    .B(_03663_),
    .X(_03765_));
 sky130_fd_sc_hd__nor2_1 _23581_ (.A(_03661_),
    .B(_03765_),
    .Y(_03766_));
 sky130_fd_sc_hd__xnor2_1 _23582_ (.A(_03764_),
    .B(_03766_),
    .Y(_03767_));
 sky130_fd_sc_hd__xnor2_1 _23583_ (.A(_03478_),
    .B(_03767_),
    .Y(_03768_));
 sky130_fd_sc_hd__xnor2_1 _23584_ (.A(_03763_),
    .B(_03768_),
    .Y(_03769_));
 sky130_fd_sc_hd__and2b_1 _23585_ (.A_N(_03666_),
    .B(_03665_),
    .X(_03770_));
 sky130_fd_sc_hd__a21oi_1 _23586_ (.A1(_03667_),
    .A2(_03672_),
    .B1(_03770_),
    .Y(_03771_));
 sky130_fd_sc_hd__xnor2_1 _23587_ (.A(_03769_),
    .B(_03771_),
    .Y(_03772_));
 sky130_fd_sc_hd__clkbuf_2 _23588_ (.A(_03583_),
    .X(_03773_));
 sky130_fd_sc_hd__nand2_1 _23589_ (.A(_03773_),
    .B(_03671_),
    .Y(_03774_));
 sky130_fd_sc_hd__a21oi_1 _23590_ (.A1(_03669_),
    .A2(_03774_),
    .B1(_03219_),
    .Y(_03775_));
 sky130_fd_sc_hd__and3_1 _23591_ (.A(_02426_),
    .B(_03669_),
    .C(_03774_),
    .X(_03776_));
 sky130_fd_sc_hd__or2_1 _23592_ (.A(_03775_),
    .B(_03776_),
    .X(_03777_));
 sky130_fd_sc_hd__xor2_1 _23593_ (.A(_03772_),
    .B(_03777_),
    .X(_03778_));
 sky130_fd_sc_hd__o21ba_1 _23594_ (.A1(_03587_),
    .A2(_03677_),
    .B1_N(_03676_),
    .X(_03779_));
 sky130_fd_sc_hd__xnor2_1 _23595_ (.A(_03778_),
    .B(_03779_),
    .Y(_03780_));
 sky130_fd_sc_hd__nand2_1 _23596_ (.A(_03585_),
    .B(_03780_),
    .Y(_03781_));
 sky130_fd_sc_hd__or2_1 _23597_ (.A(_03585_),
    .B(_03780_),
    .X(_03782_));
 sky130_fd_sc_hd__nand2_1 _23598_ (.A(_03781_),
    .B(_03782_),
    .Y(_03783_));
 sky130_fd_sc_hd__a21oi_1 _23599_ (.A1(_03680_),
    .A2(_03689_),
    .B1(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__and3_1 _23600_ (.A(_03680_),
    .B(_03689_),
    .C(_03783_),
    .X(_03785_));
 sky130_fd_sc_hd__or2_2 _23601_ (.A(_03784_),
    .B(_03785_),
    .X(_03786_));
 sky130_fd_sc_hd__o21ba_1 _23602_ (.A1(_03687_),
    .A2(_03685_),
    .B1_N(_03684_),
    .X(_03787_));
 sky130_fd_sc_hd__a21o_1 _23603_ (.A1(_03577_),
    .A2(_03686_),
    .B1(_03787_),
    .X(_03788_));
 sky130_fd_sc_hd__o31a_2 _23604_ (.A1(_03469_),
    .A2(_03470_),
    .A3(_03787_),
    .B1(_03788_),
    .X(_03789_));
 sky130_fd_sc_hd__xnor2_4 _23605_ (.A(_03786_),
    .B(_03789_),
    .Y(_00098_));
 sky130_fd_sc_hd__and2b_1 _23606_ (.A_N(_03786_),
    .B(_03789_),
    .X(_03790_));
 sky130_fd_sc_hd__or2_2 _23607_ (.A(_03784_),
    .B(_03790_),
    .X(_03791_));
 sky130_fd_sc_hd__or2b_1 _23608_ (.A(_03779_),
    .B_N(_03778_),
    .X(_03792_));
 sky130_fd_sc_hd__and2b_1 _23609_ (.A_N(_13484_),
    .B(_13803_),
    .X(_03793_));
 sky130_fd_sc_hd__nand2_1 _23610_ (.A(_13891_),
    .B(_13754_),
    .Y(_03794_));
 sky130_fd_sc_hd__xnor2_2 _23611_ (.A(_03793_),
    .B(_03794_),
    .Y(_03795_));
 sky130_fd_sc_hd__nand2_1 _23612_ (.A(_02036_),
    .B(_03695_),
    .Y(_03796_));
 sky130_fd_sc_hd__xnor2_1 _23613_ (.A(_03795_),
    .B(_03796_),
    .Y(_03797_));
 sky130_fd_sc_hd__and3_1 _23614_ (.A(_01564_),
    .B(_03287_),
    .C(_03690_),
    .X(_03798_));
 sky130_fd_sc_hd__a31o_1 _23615_ (.A1(_01885_),
    .A2(_03695_),
    .A3(_03692_),
    .B1(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__xor2_1 _23616_ (.A(_03797_),
    .B(_03799_),
    .X(_03800_));
 sky130_fd_sc_hd__a22oi_1 _23617_ (.A1(_01540_),
    .A2(_03402_),
    .B1(_03175_),
    .B2(_01544_),
    .Y(_03801_));
 sky130_fd_sc_hd__and4_1 _23618_ (.A(_14077_),
    .B(_13861_),
    .C(_13229_),
    .D(_01613_),
    .X(_03802_));
 sky130_fd_sc_hd__nor2_1 _23619_ (.A(_03801_),
    .B(_03802_),
    .Y(_03803_));
 sky130_fd_sc_hd__clkbuf_2 _23620_ (.A(_13056_),
    .X(_03804_));
 sky130_fd_sc_hd__nand2_1 _23621_ (.A(_02472_),
    .B(_03804_),
    .Y(_03805_));
 sky130_fd_sc_hd__xnor2_1 _23622_ (.A(_03803_),
    .B(_03805_),
    .Y(_03806_));
 sky130_fd_sc_hd__xnor2_1 _23623_ (.A(_03800_),
    .B(_03806_),
    .Y(_03807_));
 sky130_fd_sc_hd__and2_1 _23624_ (.A(_03694_),
    .B(_03697_),
    .X(_03808_));
 sky130_fd_sc_hd__a21oi_1 _23625_ (.A1(_03698_),
    .A2(_03703_),
    .B1(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__xor2_1 _23626_ (.A(_03807_),
    .B(_03809_),
    .X(_03810_));
 sky130_fd_sc_hd__o21ba_1 _23627_ (.A1(_03710_),
    .A2(_03713_),
    .B1_N(_03711_),
    .X(_03811_));
 sky130_fd_sc_hd__o21ba_1 _23628_ (.A1(_03699_),
    .A2(_03702_),
    .B1_N(_03700_),
    .X(_03812_));
 sky130_fd_sc_hd__a22oi_1 _23629_ (.A1(_03303_),
    .A2(_14059_),
    .B1(_01717_),
    .B2(_03503_),
    .Y(_03813_));
 sky130_fd_sc_hd__and4_1 _23630_ (.A(_03302_),
    .B(_03159_),
    .C(_01713_),
    .D(_13612_),
    .X(_03814_));
 sky130_fd_sc_hd__nor2_1 _23631_ (.A(_03813_),
    .B(_03814_),
    .Y(_03815_));
 sky130_fd_sc_hd__nand2_1 _23632_ (.A(_03307_),
    .B(_13815_),
    .Y(_03816_));
 sky130_fd_sc_hd__xnor2_1 _23633_ (.A(_03815_),
    .B(_03816_),
    .Y(_03817_));
 sky130_fd_sc_hd__xnor2_1 _23634_ (.A(_03812_),
    .B(_03817_),
    .Y(_03818_));
 sky130_fd_sc_hd__xnor2_1 _23635_ (.A(_03811_),
    .B(_03818_),
    .Y(_03819_));
 sky130_fd_sc_hd__xnor2_1 _23636_ (.A(_03810_),
    .B(_03819_),
    .Y(_03820_));
 sky130_fd_sc_hd__and2b_1 _23637_ (.A_N(_03704_),
    .B(_03706_),
    .X(_03821_));
 sky130_fd_sc_hd__a21oi_1 _23638_ (.A1(_03707_),
    .A2(_03716_),
    .B1(_03821_),
    .Y(_03822_));
 sky130_fd_sc_hd__nor2_1 _23639_ (.A(_03820_),
    .B(_03822_),
    .Y(_03823_));
 sky130_fd_sc_hd__nand2_1 _23640_ (.A(_03820_),
    .B(_03822_),
    .Y(_03824_));
 sky130_fd_sc_hd__and2b_1 _23641_ (.A_N(_03823_),
    .B(_03824_),
    .X(_03825_));
 sky130_fd_sc_hd__clkbuf_2 _23642_ (.A(_03727_),
    .X(_03826_));
 sky130_fd_sc_hd__and2b_1 _23643_ (.A_N(_03733_),
    .B(_03732_),
    .X(_03827_));
 sky130_fd_sc_hd__a21oi_1 _23644_ (.A1(_03826_),
    .A2(_03734_),
    .B1(_03827_),
    .Y(_03828_));
 sky130_fd_sc_hd__or2b_1 _23645_ (.A(_03709_),
    .B_N(_03714_),
    .X(_03829_));
 sky130_fd_sc_hd__or2b_1 _23646_ (.A(_03708_),
    .B_N(_03715_),
    .X(_03830_));
 sky130_fd_sc_hd__a22oi_2 _23647_ (.A1(_03434_),
    .A2(_13829_),
    .B1(_13831_),
    .B2(_03435_),
    .Y(_03831_));
 sky130_fd_sc_hd__and4_1 _23648_ (.A(_12324_),
    .B(_03434_),
    .C(_13826_),
    .D(_14210_),
    .X(_03832_));
 sky130_fd_sc_hd__nor2_1 _23649_ (.A(_03831_),
    .B(_03832_),
    .Y(_03833_));
 sky130_fd_sc_hd__nand2_2 _23650_ (.A(_12228_),
    .B(_14562_),
    .Y(_03834_));
 sky130_fd_sc_hd__xnor2_1 _23651_ (.A(_03833_),
    .B(_03834_),
    .Y(_03835_));
 sky130_fd_sc_hd__o21ba_1 _23652_ (.A1(_03728_),
    .A2(_03731_),
    .B1_N(_03729_),
    .X(_03836_));
 sky130_fd_sc_hd__xnor2_1 _23653_ (.A(_03835_),
    .B(_03836_),
    .Y(_03837_));
 sky130_fd_sc_hd__xnor2_1 _23654_ (.A(_03727_),
    .B(_03837_),
    .Y(_03838_));
 sky130_fd_sc_hd__a21o_1 _23655_ (.A1(_03829_),
    .A2(_03830_),
    .B1(_03838_),
    .X(_03839_));
 sky130_fd_sc_hd__nand3_1 _23656_ (.A(_03829_),
    .B(_03830_),
    .C(_03838_),
    .Y(_03840_));
 sky130_fd_sc_hd__and2_1 _23657_ (.A(_03839_),
    .B(_03840_),
    .X(_03841_));
 sky130_fd_sc_hd__xnor2_1 _23658_ (.A(_03828_),
    .B(_03841_),
    .Y(_03842_));
 sky130_fd_sc_hd__xnor2_1 _23659_ (.A(_03825_),
    .B(_03842_),
    .Y(_03843_));
 sky130_fd_sc_hd__nor2_1 _23660_ (.A(_03717_),
    .B(_03719_),
    .Y(_03844_));
 sky130_fd_sc_hd__a21oi_1 _23661_ (.A1(_03720_),
    .A2(_03739_),
    .B1(_03844_),
    .Y(_03845_));
 sky130_fd_sc_hd__xor2_1 _23662_ (.A(_03843_),
    .B(_03845_),
    .X(_03846_));
 sky130_fd_sc_hd__nor2_1 _23663_ (.A(_03238_),
    .B(_03753_),
    .Y(_03847_));
 sky130_fd_sc_hd__a21oi_1 _23664_ (.A1(_03748_),
    .A2(_03752_),
    .B1(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__or2b_1 _23665_ (.A(_03722_),
    .B_N(_03738_),
    .X(_03849_));
 sky130_fd_sc_hd__nand2_1 _23666_ (.A(_03126_),
    .B(_03377_),
    .Y(_03850_));
 sky130_fd_sc_hd__a31o_1 _23667_ (.A1(_11773_),
    .A2(_14564_),
    .A3(_03725_),
    .B1(_03629_),
    .X(_03851_));
 sky130_fd_sc_hd__nor2_1 _23668_ (.A(_03850_),
    .B(_03851_),
    .Y(_03852_));
 sky130_fd_sc_hd__o211a_1 _23669_ (.A1(_03749_),
    .A2(_03750_),
    .B1(_03851_),
    .C1(_03850_),
    .X(_03853_));
 sky130_fd_sc_hd__or2_1 _23670_ (.A(_03852_),
    .B(_03853_),
    .X(_03854_));
 sky130_fd_sc_hd__xnor2_1 _23671_ (.A(_03118_),
    .B(_03854_),
    .Y(_03855_));
 sky130_fd_sc_hd__a21oi_1 _23672_ (.A1(_03736_),
    .A2(_03849_),
    .B1(_03855_),
    .Y(_03856_));
 sky130_fd_sc_hd__and3_1 _23673_ (.A(_03736_),
    .B(_03849_),
    .C(_03855_),
    .X(_03857_));
 sky130_fd_sc_hd__nor2_1 _23674_ (.A(_03856_),
    .B(_03857_),
    .Y(_03858_));
 sky130_fd_sc_hd__xnor2_1 _23675_ (.A(_03848_),
    .B(_03858_),
    .Y(_03859_));
 sky130_fd_sc_hd__xnor2_1 _23676_ (.A(_03846_),
    .B(_03859_),
    .Y(_03860_));
 sky130_fd_sc_hd__a21oi_1 _23677_ (.A1(_03744_),
    .A2(_03756_),
    .B1(_03742_),
    .Y(_03861_));
 sky130_fd_sc_hd__nor2_1 _23678_ (.A(_03860_),
    .B(_03861_),
    .Y(_03862_));
 sky130_fd_sc_hd__and2_1 _23679_ (.A(_03860_),
    .B(_03861_),
    .X(_03863_));
 sky130_fd_sc_hd__nor2_1 _23680_ (.A(_03862_),
    .B(_03863_),
    .Y(_03864_));
 sky130_fd_sc_hd__and2b_1 _23681_ (.A_N(_03754_),
    .B(_03747_),
    .X(_03865_));
 sky130_fd_sc_hd__and2b_1 _23682_ (.A_N(_03746_),
    .B(_03755_),
    .X(_03866_));
 sky130_fd_sc_hd__nor2_1 _23683_ (.A(_03865_),
    .B(_03866_),
    .Y(_03867_));
 sky130_fd_sc_hd__xnor2_1 _23684_ (.A(_03764_),
    .B(_03867_),
    .Y(_03868_));
 sky130_fd_sc_hd__xnor2_1 _23685_ (.A(_03478_),
    .B(_03868_),
    .Y(_03869_));
 sky130_fd_sc_hd__xnor2_1 _23686_ (.A(_03864_),
    .B(_03869_),
    .Y(_03870_));
 sky130_fd_sc_hd__a21oi_1 _23687_ (.A1(_03763_),
    .A2(_03768_),
    .B1(_03761_),
    .Y(_03871_));
 sky130_fd_sc_hd__xnor2_1 _23688_ (.A(_03870_),
    .B(_03871_),
    .Y(_03872_));
 sky130_fd_sc_hd__or3_1 _23689_ (.A(_03471_),
    .B(_03472_),
    .C(_03766_),
    .X(_03873_));
 sky130_fd_sc_hd__clkbuf_2 _23690_ (.A(_03583_),
    .X(_03874_));
 sky130_fd_sc_hd__nand2_1 _23691_ (.A(_03874_),
    .B(_03767_),
    .Y(_03875_));
 sky130_fd_sc_hd__a21oi_1 _23692_ (.A1(_03873_),
    .A2(_03875_),
    .B1(_02427_),
    .Y(_03876_));
 sky130_fd_sc_hd__and3_1 _23693_ (.A(_03219_),
    .B(_03873_),
    .C(_03875_),
    .X(_03877_));
 sky130_fd_sc_hd__or2_1 _23694_ (.A(_03876_),
    .B(_03877_),
    .X(_03878_));
 sky130_fd_sc_hd__nor2_1 _23695_ (.A(_03872_),
    .B(_03878_),
    .Y(_03879_));
 sky130_fd_sc_hd__and2_1 _23696_ (.A(_03872_),
    .B(_03878_),
    .X(_03880_));
 sky130_fd_sc_hd__nor2_1 _23697_ (.A(_03879_),
    .B(_03880_),
    .Y(_03881_));
 sky130_fd_sc_hd__or2_1 _23698_ (.A(_03769_),
    .B(_03771_),
    .X(_03882_));
 sky130_fd_sc_hd__o21a_1 _23699_ (.A1(_03772_),
    .A2(_03777_),
    .B1(_03882_),
    .X(_03883_));
 sky130_fd_sc_hd__xnor2_1 _23700_ (.A(_03881_),
    .B(_03883_),
    .Y(_03884_));
 sky130_fd_sc_hd__xnor2_1 _23701_ (.A(_03775_),
    .B(_03884_),
    .Y(_03885_));
 sky130_fd_sc_hd__a21oi_1 _23702_ (.A1(_03792_),
    .A2(_03781_),
    .B1(_03885_),
    .Y(_03886_));
 sky130_fd_sc_hd__nand3_1 _23703_ (.A(_03792_),
    .B(_03781_),
    .C(_03885_),
    .Y(_03887_));
 sky130_fd_sc_hd__or2b_2 _23704_ (.A(_03886_),
    .B_N(_03887_),
    .X(_03888_));
 sky130_fd_sc_hd__xnor2_4 _23705_ (.A(_03791_),
    .B(_03888_),
    .Y(_00099_));
 sky130_fd_sc_hd__or3_1 _23706_ (.A(_03879_),
    .B(_03880_),
    .C(_03883_),
    .X(_03889_));
 sky130_fd_sc_hd__nand2_1 _23707_ (.A(_03775_),
    .B(_03884_),
    .Y(_03890_));
 sky130_fd_sc_hd__and2b_1 _23708_ (.A_N(_14268_),
    .B(_13803_),
    .X(_03891_));
 sky130_fd_sc_hd__a21oi_1 _23709_ (.A1(_14081_),
    .A2(_13754_),
    .B1(_03891_),
    .Y(_03892_));
 sky130_fd_sc_hd__and3_1 _23710_ (.A(_14444_),
    .B(_01625_),
    .C(_03891_),
    .X(_03893_));
 sky130_fd_sc_hd__nor2_1 _23711_ (.A(_03892_),
    .B(_03893_),
    .Y(_03894_));
 sky130_fd_sc_hd__nand2_1 _23712_ (.A(_03308_),
    .B(_03286_),
    .Y(_03895_));
 sky130_fd_sc_hd__xnor2_2 _23713_ (.A(_03894_),
    .B(_03895_),
    .Y(_03896_));
 sky130_fd_sc_hd__and3_1 _23714_ (.A(_01885_),
    .B(_03287_),
    .C(_03793_),
    .X(_03897_));
 sky130_fd_sc_hd__a31oi_4 _23715_ (.A1(_02036_),
    .A2(_03695_),
    .A3(_03795_),
    .B1(_03897_),
    .Y(_03898_));
 sky130_fd_sc_hd__xnor2_2 _23716_ (.A(_03896_),
    .B(_03898_),
    .Y(_03899_));
 sky130_fd_sc_hd__a22oi_1 _23717_ (.A1(_01538_),
    .A2(_03402_),
    .B1(_03175_),
    .B2(_01540_),
    .Y(_03900_));
 sky130_fd_sc_hd__and4_1 _23718_ (.A(_13864_),
    .B(_13868_),
    .C(_13224_),
    .D(_14510_),
    .X(_03901_));
 sky130_fd_sc_hd__or2_1 _23719_ (.A(_03900_),
    .B(_03901_),
    .X(_03902_));
 sky130_fd_sc_hd__nand2_1 _23720_ (.A(_03179_),
    .B(_02610_),
    .Y(_03903_));
 sky130_fd_sc_hd__xor2_2 _23721_ (.A(_03902_),
    .B(_03903_),
    .X(_03904_));
 sky130_fd_sc_hd__xnor2_2 _23722_ (.A(_03899_),
    .B(_03904_),
    .Y(_03905_));
 sky130_fd_sc_hd__and2_1 _23723_ (.A(_03797_),
    .B(_03799_),
    .X(_03906_));
 sky130_fd_sc_hd__a21oi_2 _23724_ (.A1(_03800_),
    .A2(_03806_),
    .B1(_03906_),
    .Y(_03907_));
 sky130_fd_sc_hd__xor2_1 _23725_ (.A(_03905_),
    .B(_03907_),
    .X(_03908_));
 sky130_fd_sc_hd__a31o_1 _23726_ (.A1(_12587_),
    .A2(_13816_),
    .A3(_03815_),
    .B1(_03814_),
    .X(_03909_));
 sky130_fd_sc_hd__a31o_1 _23727_ (.A1(_02472_),
    .A2(_03804_),
    .A3(_03803_),
    .B1(_03802_),
    .X(_03910_));
 sky130_fd_sc_hd__a22oi_1 _23728_ (.A1(_03303_),
    .A2(_01717_),
    .B1(_01870_),
    .B2(_03503_),
    .Y(_03911_));
 sky130_fd_sc_hd__and4_1 _23729_ (.A(_12772_),
    .B(_13961_),
    .C(_13836_),
    .D(_13824_),
    .X(_03912_));
 sky130_fd_sc_hd__nor2_1 _23730_ (.A(_03911_),
    .B(_03912_),
    .Y(_03913_));
 sky130_fd_sc_hd__nand2_1 _23731_ (.A(_03307_),
    .B(_14023_),
    .Y(_03914_));
 sky130_fd_sc_hd__xnor2_1 _23732_ (.A(_03913_),
    .B(_03914_),
    .Y(_03915_));
 sky130_fd_sc_hd__xor2_1 _23733_ (.A(_03910_),
    .B(_03915_),
    .X(_03916_));
 sky130_fd_sc_hd__nand2_1 _23734_ (.A(_03909_),
    .B(_03916_),
    .Y(_03917_));
 sky130_fd_sc_hd__or2_1 _23735_ (.A(_03909_),
    .B(_03916_),
    .X(_03918_));
 sky130_fd_sc_hd__and2_1 _23736_ (.A(_03917_),
    .B(_03918_),
    .X(_03919_));
 sky130_fd_sc_hd__xnor2_1 _23737_ (.A(_03908_),
    .B(_03919_),
    .Y(_03920_));
 sky130_fd_sc_hd__nor2_1 _23738_ (.A(_03807_),
    .B(_03809_),
    .Y(_03921_));
 sky130_fd_sc_hd__a21oi_2 _23739_ (.A1(_03810_),
    .A2(_03819_),
    .B1(_03921_),
    .Y(_03922_));
 sky130_fd_sc_hd__xor2_1 _23740_ (.A(_03920_),
    .B(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__or2b_1 _23741_ (.A(_03836_),
    .B_N(_03835_),
    .X(_03924_));
 sky130_fd_sc_hd__a21bo_1 _23742_ (.A1(_03826_),
    .A2(_03837_),
    .B1_N(_03924_),
    .X(_03925_));
 sky130_fd_sc_hd__or2b_1 _23743_ (.A(_03812_),
    .B_N(_03817_),
    .X(_03926_));
 sky130_fd_sc_hd__or2b_1 _23744_ (.A(_03811_),
    .B_N(_03818_),
    .X(_03927_));
 sky130_fd_sc_hd__nand2_1 _23745_ (.A(_03926_),
    .B(_03927_),
    .Y(_03928_));
 sky130_fd_sc_hd__o21ba_1 _23746_ (.A1(_03831_),
    .A2(_03834_),
    .B1_N(_03832_),
    .X(_03929_));
 sky130_fd_sc_hd__a22o_1 _23747_ (.A1(_03633_),
    .A2(_14211_),
    .B1(_14037_),
    .B2(_03435_),
    .X(_03930_));
 sky130_fd_sc_hd__nand4_1 _23748_ (.A(_12325_),
    .B(_03633_),
    .C(_03547_),
    .D(_14562_),
    .Y(_03931_));
 sky130_fd_sc_hd__nand2_1 _23749_ (.A(_03930_),
    .B(_03931_),
    .Y(_03932_));
 sky130_fd_sc_hd__xor2_1 _23750_ (.A(_03834_),
    .B(_03932_),
    .X(_03933_));
 sky130_fd_sc_hd__xnor2_1 _23751_ (.A(_03929_),
    .B(_03933_),
    .Y(_03934_));
 sky130_fd_sc_hd__xnor2_1 _23752_ (.A(_03727_),
    .B(_03934_),
    .Y(_03935_));
 sky130_fd_sc_hd__xnor2_1 _23753_ (.A(_03928_),
    .B(_03935_),
    .Y(_03936_));
 sky130_fd_sc_hd__xnor2_1 _23754_ (.A(_03925_),
    .B(_03936_),
    .Y(_03937_));
 sky130_vsdinv _23755_ (.A(_03937_),
    .Y(_03938_));
 sky130_fd_sc_hd__xnor2_1 _23756_ (.A(_03923_),
    .B(_03938_),
    .Y(_03939_));
 sky130_fd_sc_hd__a21oi_1 _23757_ (.A1(_03824_),
    .A2(_03842_),
    .B1(_03823_),
    .Y(_03940_));
 sky130_fd_sc_hd__nor2_1 _23758_ (.A(_03939_),
    .B(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__and2_1 _23759_ (.A(_03939_),
    .B(_03940_),
    .X(_03942_));
 sky130_fd_sc_hd__or2_1 _23760_ (.A(_03941_),
    .B(_03942_),
    .X(_03943_));
 sky130_fd_sc_hd__nand2_1 _23761_ (.A(_03750_),
    .B(_03851_),
    .Y(_03944_));
 sky130_fd_sc_hd__o21ai_1 _23762_ (.A1(_03238_),
    .A2(_03854_),
    .B1(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__or2b_1 _23763_ (.A(_03828_),
    .B_N(_03841_),
    .X(_03946_));
 sky130_fd_sc_hd__nand2_1 _23764_ (.A(_03839_),
    .B(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__and2_1 _23765_ (.A(_03750_),
    .B(_03851_),
    .X(_03948_));
 sky130_fd_sc_hd__or2_1 _23766_ (.A(_03852_),
    .B(_03948_),
    .X(_03949_));
 sky130_fd_sc_hd__xnor2_2 _23767_ (.A(_03118_),
    .B(_03949_),
    .Y(_03950_));
 sky130_fd_sc_hd__xnor2_1 _23768_ (.A(_03947_),
    .B(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__xnor2_1 _23769_ (.A(_03945_),
    .B(_03951_),
    .Y(_03952_));
 sky130_fd_sc_hd__xnor2_1 _23770_ (.A(_03943_),
    .B(_03952_),
    .Y(_03953_));
 sky130_fd_sc_hd__nor2_1 _23771_ (.A(_03843_),
    .B(_03845_),
    .Y(_03954_));
 sky130_fd_sc_hd__a21oi_1 _23772_ (.A1(_03846_),
    .A2(_03859_),
    .B1(_03954_),
    .Y(_03955_));
 sky130_fd_sc_hd__xor2_1 _23773_ (.A(_03953_),
    .B(_03955_),
    .X(_03956_));
 sky130_fd_sc_hd__and2b_1 _23774_ (.A_N(_03848_),
    .B(_03858_),
    .X(_03957_));
 sky130_fd_sc_hd__nor2_1 _23775_ (.A(_03856_),
    .B(_03957_),
    .Y(_03958_));
 sky130_fd_sc_hd__xnor2_1 _23776_ (.A(_03368_),
    .B(_03958_),
    .Y(_03959_));
 sky130_fd_sc_hd__xnor2_1 _23777_ (.A(_03478_),
    .B(_03959_),
    .Y(_03960_));
 sky130_fd_sc_hd__xnor2_1 _23778_ (.A(_03956_),
    .B(_03960_),
    .Y(_03961_));
 sky130_fd_sc_hd__a21oi_1 _23779_ (.A1(_03864_),
    .A2(_03869_),
    .B1(_03862_),
    .Y(_03962_));
 sky130_fd_sc_hd__xnor2_1 _23780_ (.A(_03961_),
    .B(_03962_),
    .Y(_03963_));
 sky130_fd_sc_hd__or3_1 _23781_ (.A(_03471_),
    .B(_03472_),
    .C(_03867_),
    .X(_03964_));
 sky130_fd_sc_hd__nand2_1 _23782_ (.A(_03773_),
    .B(_03868_),
    .Y(_03965_));
 sky130_fd_sc_hd__a21oi_1 _23783_ (.A1(_03964_),
    .A2(_03965_),
    .B1(_03219_),
    .Y(_03966_));
 sky130_fd_sc_hd__and3_1 _23784_ (.A(_02426_),
    .B(_03964_),
    .C(_03965_),
    .X(_03967_));
 sky130_fd_sc_hd__or2_1 _23785_ (.A(_03966_),
    .B(_03967_),
    .X(_03968_));
 sky130_fd_sc_hd__nor2_1 _23786_ (.A(_03963_),
    .B(_03968_),
    .Y(_03969_));
 sky130_fd_sc_hd__and2_1 _23787_ (.A(_03963_),
    .B(_03968_),
    .X(_03970_));
 sky130_fd_sc_hd__nor2_1 _23788_ (.A(_03969_),
    .B(_03970_),
    .Y(_03971_));
 sky130_fd_sc_hd__o21ba_1 _23789_ (.A1(_03870_),
    .A2(_03871_),
    .B1_N(_03879_),
    .X(_03972_));
 sky130_fd_sc_hd__xnor2_1 _23790_ (.A(_03971_),
    .B(_03972_),
    .Y(_03973_));
 sky130_fd_sc_hd__nand2_1 _23791_ (.A(_03876_),
    .B(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__or2_1 _23792_ (.A(_03876_),
    .B(_03973_),
    .X(_03975_));
 sky130_fd_sc_hd__nand2_1 _23793_ (.A(_03974_),
    .B(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__a21o_1 _23794_ (.A1(_03889_),
    .A2(_03890_),
    .B1(_03976_),
    .X(_03977_));
 sky130_fd_sc_hd__and3_1 _23795_ (.A(_03889_),
    .B(_03890_),
    .C(_03976_),
    .X(_03978_));
 sky130_vsdinv _23796_ (.A(_03978_),
    .Y(_03979_));
 sky130_fd_sc_hd__nand2_2 _23797_ (.A(_03977_),
    .B(_03979_),
    .Y(_03980_));
 sky130_fd_sc_hd__nor2_1 _23798_ (.A(_03786_),
    .B(_03888_),
    .Y(_03981_));
 sky130_fd_sc_hd__o311ai_4 _23799_ (.A1(_03469_),
    .A2(_03470_),
    .A3(_03787_),
    .B1(_03788_),
    .C1(_03981_),
    .Y(_03982_));
 sky130_fd_sc_hd__o21ai_1 _23800_ (.A1(_03784_),
    .A2(_03886_),
    .B1(_03887_),
    .Y(_03983_));
 sky130_fd_sc_hd__nand2_2 _23801_ (.A(_03982_),
    .B(_03983_),
    .Y(_03984_));
 sky130_fd_sc_hd__xnor2_4 _23802_ (.A(_03980_),
    .B(_03984_),
    .Y(_00100_));
 sky130_fd_sc_hd__or3_1 _23803_ (.A(_03969_),
    .B(_03970_),
    .C(_03972_),
    .X(_03985_));
 sky130_fd_sc_hd__and2b_1 _23804_ (.A_N(_14080_),
    .B(_13803_),
    .X(_03986_));
 sky130_fd_sc_hd__a21oi_1 _23805_ (.A1(_03308_),
    .A2(_03287_),
    .B1(_03986_),
    .Y(_03987_));
 sky130_fd_sc_hd__and3_1 _23806_ (.A(_14077_),
    .B(_03287_),
    .C(_03986_),
    .X(_03988_));
 sky130_fd_sc_hd__nor2_1 _23807_ (.A(_03987_),
    .B(_03988_),
    .Y(_03989_));
 sky130_fd_sc_hd__nand2_1 _23808_ (.A(_02331_),
    .B(_03695_),
    .Y(_03990_));
 sky130_fd_sc_hd__xnor2_1 _23809_ (.A(_03989_),
    .B(_03990_),
    .Y(_03991_));
 sky130_fd_sc_hd__o21ba_1 _23810_ (.A1(_03892_),
    .A2(_03895_),
    .B1_N(_03893_),
    .X(_03992_));
 sky130_fd_sc_hd__xnor2_1 _23811_ (.A(_03991_),
    .B(_03992_),
    .Y(_03993_));
 sky130_fd_sc_hd__a22oi_1 _23812_ (.A1(_02610_),
    .A2(_03596_),
    .B1(_03597_),
    .B2(_13869_),
    .Y(_03994_));
 sky130_fd_sc_hd__and4_1 _23813_ (.A(_14438_),
    .B(_01866_),
    .C(_03402_),
    .D(_03175_),
    .X(_03995_));
 sky130_fd_sc_hd__or2_1 _23814_ (.A(_03994_),
    .B(_03995_),
    .X(_03996_));
 sky130_fd_sc_hd__nand2_1 _23815_ (.A(_03804_),
    .B(_01718_),
    .Y(_03997_));
 sky130_fd_sc_hd__xor2_1 _23816_ (.A(_03996_),
    .B(_03997_),
    .X(_03998_));
 sky130_fd_sc_hd__xnor2_1 _23817_ (.A(_03993_),
    .B(_03998_),
    .Y(_03999_));
 sky130_fd_sc_hd__and2b_1 _23818_ (.A_N(_03898_),
    .B(_03896_),
    .X(_04000_));
 sky130_fd_sc_hd__a21oi_1 _23819_ (.A1(_03899_),
    .A2(_03904_),
    .B1(_04000_),
    .Y(_04001_));
 sky130_fd_sc_hd__nor2_1 _23820_ (.A(_03999_),
    .B(_04001_),
    .Y(_04002_));
 sky130_fd_sc_hd__nand2_1 _23821_ (.A(_03999_),
    .B(_04001_),
    .Y(_04003_));
 sky130_fd_sc_hd__and2b_1 _23822_ (.A_N(_04002_),
    .B(_04003_),
    .X(_04004_));
 sky130_fd_sc_hd__a31o_1 _23823_ (.A1(_12587_),
    .A2(_13819_),
    .A3(_03913_),
    .B1(_03912_),
    .X(_04005_));
 sky130_fd_sc_hd__nor2_1 _23824_ (.A(_03902_),
    .B(_03903_),
    .Y(_04006_));
 sky130_fd_sc_hd__a22oi_1 _23825_ (.A1(_03159_),
    .A2(_01870_),
    .B1(_13829_),
    .B2(_03302_),
    .Y(_04007_));
 sky130_fd_sc_hd__and4_1 _23826_ (.A(_12772_),
    .B(_13961_),
    .C(_13824_),
    .D(_01846_),
    .X(_04008_));
 sky130_fd_sc_hd__o2bb2a_1 _23827_ (.A1_N(_12586_),
    .A2_N(_03547_),
    .B1(_04007_),
    .B2(_04008_),
    .X(_04009_));
 sky130_fd_sc_hd__and4bb_1 _23828_ (.A_N(_04007_),
    .B_N(_04008_),
    .C(_12586_),
    .D(_14211_),
    .X(_04010_));
 sky130_fd_sc_hd__nor2_1 _23829_ (.A(_04009_),
    .B(_04010_),
    .Y(_04011_));
 sky130_fd_sc_hd__o21ai_2 _23830_ (.A1(_03901_),
    .A2(_04006_),
    .B1(_04011_),
    .Y(_04012_));
 sky130_fd_sc_hd__or3_1 _23831_ (.A(_03901_),
    .B(_04006_),
    .C(_04011_),
    .X(_04013_));
 sky130_fd_sc_hd__and2_1 _23832_ (.A(_04012_),
    .B(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__nand2_1 _23833_ (.A(_04005_),
    .B(_04014_),
    .Y(_04015_));
 sky130_fd_sc_hd__or2_1 _23834_ (.A(_04005_),
    .B(_04014_),
    .X(_04016_));
 sky130_fd_sc_hd__and2_1 _23835_ (.A(_04015_),
    .B(_04016_),
    .X(_04017_));
 sky130_fd_sc_hd__xnor2_2 _23836_ (.A(_04004_),
    .B(_04017_),
    .Y(_04018_));
 sky130_fd_sc_hd__nor2_1 _23837_ (.A(_03905_),
    .B(_03907_),
    .Y(_04019_));
 sky130_fd_sc_hd__a21oi_1 _23838_ (.A1(_03908_),
    .A2(_03919_),
    .B1(_04019_),
    .Y(_04020_));
 sky130_fd_sc_hd__xnor2_1 _23839_ (.A(_04018_),
    .B(_04020_),
    .Y(_04021_));
 sky130_fd_sc_hd__and2b_1 _23840_ (.A_N(_03929_),
    .B(_03933_),
    .X(_04022_));
 sky130_fd_sc_hd__a21oi_1 _23841_ (.A1(_03826_),
    .A2(_03934_),
    .B1(_04022_),
    .Y(_04023_));
 sky130_fd_sc_hd__nand2_1 _23842_ (.A(_03910_),
    .B(_03915_),
    .Y(_04024_));
 sky130_fd_sc_hd__and3_1 _23843_ (.A(_12325_),
    .B(_03633_),
    .C(_14563_),
    .X(_04025_));
 sky130_fd_sc_hd__o21ai_1 _23844_ (.A1(_12325_),
    .A2(_03633_),
    .B1(_14563_),
    .Y(_04026_));
 sky130_fd_sc_hd__nor2_1 _23845_ (.A(_04025_),
    .B(_04026_),
    .Y(_04027_));
 sky130_fd_sc_hd__o22a_1 _23846_ (.A1(_03834_),
    .A2(_03930_),
    .B1(_03931_),
    .B2(_12229_),
    .X(_04028_));
 sky130_fd_sc_hd__xnor2_1 _23847_ (.A(_04027_),
    .B(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__xnor2_1 _23848_ (.A(_03727_),
    .B(_04029_),
    .Y(_04030_));
 sky130_fd_sc_hd__a21oi_1 _23849_ (.A1(_04024_),
    .A2(_03917_),
    .B1(_04030_),
    .Y(_04031_));
 sky130_fd_sc_hd__and3_1 _23850_ (.A(_04024_),
    .B(_03917_),
    .C(_04030_),
    .X(_04032_));
 sky130_fd_sc_hd__nor2_1 _23851_ (.A(_04031_),
    .B(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__xnor2_1 _23852_ (.A(_04023_),
    .B(_04033_),
    .Y(_04034_));
 sky130_fd_sc_hd__xnor2_1 _23853_ (.A(_04021_),
    .B(_04034_),
    .Y(_04035_));
 sky130_fd_sc_hd__nor2_1 _23854_ (.A(_03920_),
    .B(_03922_),
    .Y(_04036_));
 sky130_fd_sc_hd__a21oi_1 _23855_ (.A1(_03923_),
    .A2(_03938_),
    .B1(_04036_),
    .Y(_04037_));
 sky130_fd_sc_hd__xor2_1 _23856_ (.A(_04035_),
    .B(_04037_),
    .X(_04038_));
 sky130_fd_sc_hd__o21a_1 _23857_ (.A1(_03238_),
    .A2(_03852_),
    .B1(_03944_),
    .X(_04039_));
 sky130_fd_sc_hd__clkbuf_2 _23858_ (.A(_04039_),
    .X(_04040_));
 sky130_fd_sc_hd__a21oi_1 _23859_ (.A1(_03926_),
    .A2(_03927_),
    .B1(_03935_),
    .Y(_04041_));
 sky130_fd_sc_hd__a21oi_1 _23860_ (.A1(_03925_),
    .A2(_03936_),
    .B1(_04041_),
    .Y(_04042_));
 sky130_fd_sc_hd__or2_1 _23861_ (.A(_03950_),
    .B(_04042_),
    .X(_04043_));
 sky130_fd_sc_hd__clkbuf_2 _23862_ (.A(_03950_),
    .X(_04044_));
 sky130_fd_sc_hd__nand2_1 _23863_ (.A(_04044_),
    .B(_04042_),
    .Y(_04045_));
 sky130_fd_sc_hd__nand2_1 _23864_ (.A(_04043_),
    .B(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hd__xor2_1 _23865_ (.A(_04040_),
    .B(_04046_),
    .X(_04047_));
 sky130_fd_sc_hd__xnor2_1 _23866_ (.A(_04038_),
    .B(_04047_),
    .Y(_04048_));
 sky130_fd_sc_hd__o21ba_1 _23867_ (.A1(_03943_),
    .A2(_03952_),
    .B1_N(_03941_),
    .X(_04049_));
 sky130_fd_sc_hd__xnor2_1 _23868_ (.A(_04048_),
    .B(_04049_),
    .Y(_04050_));
 sky130_fd_sc_hd__a21oi_1 _23869_ (.A1(_03839_),
    .A2(_03946_),
    .B1(_04044_),
    .Y(_04051_));
 sky130_fd_sc_hd__a21o_1 _23870_ (.A1(_03945_),
    .A2(_03951_),
    .B1(_04051_),
    .X(_04052_));
 sky130_fd_sc_hd__xor2_1 _23871_ (.A(_03368_),
    .B(_04052_),
    .X(_04053_));
 sky130_fd_sc_hd__nand2_1 _23872_ (.A(_03583_),
    .B(_04053_),
    .Y(_04054_));
 sky130_fd_sc_hd__or2_1 _23873_ (.A(_03583_),
    .B(_04053_),
    .X(_04055_));
 sky130_fd_sc_hd__and2_1 _23874_ (.A(_04054_),
    .B(_04055_),
    .X(_04056_));
 sky130_fd_sc_hd__xnor2_1 _23875_ (.A(_04050_),
    .B(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__nor2_1 _23876_ (.A(_03953_),
    .B(_03955_),
    .Y(_04058_));
 sky130_fd_sc_hd__a21oi_1 _23877_ (.A1(_03956_),
    .A2(_03960_),
    .B1(_04058_),
    .Y(_04059_));
 sky130_fd_sc_hd__xnor2_1 _23878_ (.A(_04057_),
    .B(_04059_),
    .Y(_04060_));
 sky130_fd_sc_hd__or3_1 _23879_ (.A(_03471_),
    .B(_03472_),
    .C(_03958_),
    .X(_04061_));
 sky130_fd_sc_hd__nand2_1 _23880_ (.A(_03773_),
    .B(_03959_),
    .Y(_04062_));
 sky130_fd_sc_hd__a21oi_1 _23881_ (.A1(_04061_),
    .A2(_04062_),
    .B1(_03219_),
    .Y(_04063_));
 sky130_fd_sc_hd__and3_1 _23882_ (.A(_02426_),
    .B(_04061_),
    .C(_04062_),
    .X(_04064_));
 sky130_fd_sc_hd__or2_1 _23883_ (.A(_04063_),
    .B(_04064_),
    .X(_04065_));
 sky130_fd_sc_hd__nor2_1 _23884_ (.A(_04060_),
    .B(_04065_),
    .Y(_04066_));
 sky130_fd_sc_hd__and2_1 _23885_ (.A(_04060_),
    .B(_04065_),
    .X(_04067_));
 sky130_fd_sc_hd__nor2_1 _23886_ (.A(_04066_),
    .B(_04067_),
    .Y(_04068_));
 sky130_fd_sc_hd__o21ba_1 _23887_ (.A1(_03961_),
    .A2(_03962_),
    .B1_N(_03969_),
    .X(_04069_));
 sky130_fd_sc_hd__xnor2_1 _23888_ (.A(_04068_),
    .B(_04069_),
    .Y(_04070_));
 sky130_fd_sc_hd__nand2_1 _23889_ (.A(_03966_),
    .B(_04070_),
    .Y(_04071_));
 sky130_fd_sc_hd__or2_1 _23890_ (.A(_03966_),
    .B(_04070_),
    .X(_04072_));
 sky130_fd_sc_hd__nand2_1 _23891_ (.A(_04071_),
    .B(_04072_),
    .Y(_04073_));
 sky130_fd_sc_hd__and3_1 _23892_ (.A(_03985_),
    .B(_03974_),
    .C(_04073_),
    .X(_04074_));
 sky130_fd_sc_hd__a21o_1 _23893_ (.A1(_03985_),
    .A2(_03974_),
    .B1(_04073_),
    .X(_04075_));
 sky130_fd_sc_hd__or2b_2 _23894_ (.A(_04074_),
    .B_N(_04075_),
    .X(_04076_));
 sky130_fd_sc_hd__a21bo_1 _23895_ (.A1(_03979_),
    .A2(_03984_),
    .B1_N(_03977_),
    .X(_04077_));
 sky130_fd_sc_hd__xnor2_4 _23896_ (.A(_04076_),
    .B(_04077_),
    .Y(_00101_));
 sky130_fd_sc_hd__or3_1 _23897_ (.A(_04066_),
    .B(_04067_),
    .C(_04069_),
    .X(_04078_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _23898_ (.A(_01625_),
    .X(_04079_));
 sky130_fd_sc_hd__and2b_1 _23899_ (.A_N(_01544_),
    .B(_13804_),
    .X(_04080_));
 sky130_fd_sc_hd__a21oi_1 _23900_ (.A1(_02331_),
    .A2(_04079_),
    .B1(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__and3_1 _23901_ (.A(_02331_),
    .B(_04079_),
    .C(_04080_),
    .X(_04082_));
 sky130_fd_sc_hd__nor2_1 _23902_ (.A(_04081_),
    .B(_04082_),
    .Y(_04083_));
 sky130_fd_sc_hd__clkbuf_2 _23903_ (.A(_03695_),
    .X(_04084_));
 sky130_fd_sc_hd__nand2_1 _23904_ (.A(_02472_),
    .B(_04084_),
    .Y(_04085_));
 sky130_fd_sc_hd__xnor2_1 _23905_ (.A(_04083_),
    .B(_04085_),
    .Y(_04086_));
 sky130_fd_sc_hd__o21ba_1 _23906_ (.A1(_03987_),
    .A2(_03990_),
    .B1_N(_03988_),
    .X(_04087_));
 sky130_fd_sc_hd__xnor2_1 _23907_ (.A(_04086_),
    .B(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hd__buf_2 _23908_ (.A(_03596_),
    .X(_04089_));
 sky130_fd_sc_hd__clkbuf_2 _23909_ (.A(_01844_),
    .X(_04090_));
 sky130_fd_sc_hd__clkbuf_4 _23910_ (.A(_03597_),
    .X(_04091_));
 sky130_fd_sc_hd__clkbuf_2 _23911_ (.A(_02610_),
    .X(_04092_));
 sky130_fd_sc_hd__a22oi_1 _23912_ (.A1(_04089_),
    .A2(_04090_),
    .B1(_04091_),
    .B2(_04092_),
    .Y(_04093_));
 sky130_fd_sc_hd__buf_1 _23913_ (.A(_03596_),
    .X(_04094_));
 sky130_fd_sc_hd__buf_1 _23914_ (.A(_03597_),
    .X(_04095_));
 sky130_fd_sc_hd__and4_1 _23915_ (.A(_04092_),
    .B(_04094_),
    .C(_04090_),
    .D(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__nor2_1 _23916_ (.A(_04093_),
    .B(_04096_),
    .Y(_04097_));
 sky130_fd_sc_hd__clkbuf_4 _23917_ (.A(_03804_),
    .X(_04098_));
 sky130_fd_sc_hd__nand2_1 _23918_ (.A(_04098_),
    .B(_13816_),
    .Y(_04099_));
 sky130_fd_sc_hd__xnor2_1 _23919_ (.A(_04097_),
    .B(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__xnor2_1 _23920_ (.A(_04088_),
    .B(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__and2b_1 _23921_ (.A_N(_03992_),
    .B(_03991_),
    .X(_04102_));
 sky130_fd_sc_hd__a21oi_1 _23922_ (.A1(_03993_),
    .A2(_03998_),
    .B1(_04102_),
    .Y(_04103_));
 sky130_fd_sc_hd__xor2_1 _23923_ (.A(_04101_),
    .B(_04103_),
    .X(_04104_));
 sky130_fd_sc_hd__nor2_1 _23924_ (.A(_03996_),
    .B(_03997_),
    .Y(_04105_));
 sky130_fd_sc_hd__a22oi_1 _23925_ (.A1(_03609_),
    .A2(_13817_),
    .B1(_14211_),
    .B2(_12773_),
    .Y(_04106_));
 sky130_fd_sc_hd__and4_1 _23926_ (.A(_03503_),
    .B(_03303_),
    .C(_13829_),
    .D(_13827_),
    .X(_04107_));
 sky130_fd_sc_hd__nor2_1 _23927_ (.A(_04106_),
    .B(_04107_),
    .Y(_04108_));
 sky130_fd_sc_hd__nand2_4 _23928_ (.A(_03307_),
    .B(_14562_),
    .Y(_04109_));
 sky130_fd_sc_hd__xnor2_1 _23929_ (.A(_04108_),
    .B(_04109_),
    .Y(_04110_));
 sky130_fd_sc_hd__o21ai_2 _23930_ (.A1(_03995_),
    .A2(_04105_),
    .B1(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__or3_1 _23931_ (.A(_03995_),
    .B(_04105_),
    .C(_04110_),
    .X(_04112_));
 sky130_fd_sc_hd__and2_1 _23932_ (.A(_04111_),
    .B(_04112_),
    .X(_04113_));
 sky130_fd_sc_hd__o21ai_1 _23933_ (.A1(_04008_),
    .A2(_04010_),
    .B1(_04113_),
    .Y(_04114_));
 sky130_fd_sc_hd__or3_1 _23934_ (.A(_04008_),
    .B(_04010_),
    .C(_04113_),
    .X(_04115_));
 sky130_fd_sc_hd__and2_1 _23935_ (.A(_04114_),
    .B(_04115_),
    .X(_04116_));
 sky130_fd_sc_hd__xnor2_1 _23936_ (.A(_04104_),
    .B(_04116_),
    .Y(_04117_));
 sky130_fd_sc_hd__a21oi_2 _23937_ (.A1(_04003_),
    .A2(_04017_),
    .B1(_04002_),
    .Y(_04118_));
 sky130_fd_sc_hd__xor2_1 _23938_ (.A(_04117_),
    .B(_04118_),
    .X(_04119_));
 sky130_fd_sc_hd__and2_1 _23939_ (.A(_12229_),
    .B(_04025_),
    .X(_04120_));
 sky130_fd_sc_hd__a21oi_1 _23940_ (.A1(_03826_),
    .A2(_04029_),
    .B1(_04120_),
    .Y(_04121_));
 sky130_fd_sc_hd__nand2_1 _23941_ (.A(_03834_),
    .B(_04026_),
    .Y(_04122_));
 sky130_fd_sc_hd__and2b_1 _23942_ (.A_N(_04120_),
    .B(_04122_),
    .X(_04123_));
 sky130_fd_sc_hd__xnor2_2 _23943_ (.A(_03826_),
    .B(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hd__a21oi_1 _23944_ (.A1(_04012_),
    .A2(_04015_),
    .B1(_04124_),
    .Y(_04125_));
 sky130_fd_sc_hd__and3_1 _23945_ (.A(_04012_),
    .B(_04015_),
    .C(_04124_),
    .X(_04126_));
 sky130_fd_sc_hd__nor2_1 _23946_ (.A(_04125_),
    .B(_04126_),
    .Y(_04127_));
 sky130_fd_sc_hd__xnor2_1 _23947_ (.A(_04121_),
    .B(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hd__xnor2_1 _23948_ (.A(_04119_),
    .B(_04128_),
    .Y(_04129_));
 sky130_fd_sc_hd__nand2_1 _23949_ (.A(_04018_),
    .B(_04020_),
    .Y(_04130_));
 sky130_fd_sc_hd__nor2_1 _23950_ (.A(_04018_),
    .B(_04020_),
    .Y(_04131_));
 sky130_fd_sc_hd__a21oi_1 _23951_ (.A1(_04130_),
    .A2(_04034_),
    .B1(_04131_),
    .Y(_04132_));
 sky130_fd_sc_hd__xor2_1 _23952_ (.A(_04129_),
    .B(_04132_),
    .X(_04133_));
 sky130_fd_sc_hd__and2b_1 _23953_ (.A_N(_04023_),
    .B(_04033_),
    .X(_04134_));
 sky130_fd_sc_hd__nor2_1 _23954_ (.A(_04031_),
    .B(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__xnor2_1 _23955_ (.A(_03950_),
    .B(_04135_),
    .Y(_04136_));
 sky130_fd_sc_hd__or2_1 _23956_ (.A(_04039_),
    .B(_04136_),
    .X(_04137_));
 sky130_fd_sc_hd__nand2_1 _23957_ (.A(_04040_),
    .B(_04136_),
    .Y(_04138_));
 sky130_fd_sc_hd__and2_1 _23958_ (.A(_04137_),
    .B(_04138_),
    .X(_04139_));
 sky130_fd_sc_hd__xnor2_1 _23959_ (.A(_04133_),
    .B(_04139_),
    .Y(_04140_));
 sky130_fd_sc_hd__or2b_1 _23960_ (.A(_04035_),
    .B_N(_04037_),
    .X(_04141_));
 sky130_fd_sc_hd__and2b_1 _23961_ (.A_N(_04037_),
    .B(_04035_),
    .X(_04142_));
 sky130_fd_sc_hd__a21oi_1 _23962_ (.A1(_04141_),
    .A2(_04047_),
    .B1(_04142_),
    .Y(_04143_));
 sky130_fd_sc_hd__xor2_1 _23963_ (.A(_04140_),
    .B(_04143_),
    .X(_04144_));
 sky130_fd_sc_hd__o21a_1 _23964_ (.A1(_04040_),
    .A2(_04046_),
    .B1(_04043_),
    .X(_04145_));
 sky130_fd_sc_hd__xnor2_1 _23965_ (.A(_03764_),
    .B(_04145_),
    .Y(_04146_));
 sky130_fd_sc_hd__nand2_1 _23966_ (.A(_03773_),
    .B(_04146_),
    .Y(_04147_));
 sky130_fd_sc_hd__or2_1 _23967_ (.A(_03583_),
    .B(_04146_),
    .X(_04148_));
 sky130_fd_sc_hd__and2_1 _23968_ (.A(_04147_),
    .B(_04148_),
    .X(_04149_));
 sky130_fd_sc_hd__xnor2_1 _23969_ (.A(_04144_),
    .B(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hd__and2b_1 _23970_ (.A_N(_04049_),
    .B(_04048_),
    .X(_04151_));
 sky130_fd_sc_hd__a21oi_1 _23971_ (.A1(_04050_),
    .A2(_04056_),
    .B1(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__or2_1 _23972_ (.A(_04150_),
    .B(_04152_),
    .X(_04153_));
 sky130_fd_sc_hd__nand2_1 _23973_ (.A(_04150_),
    .B(_04152_),
    .Y(_04154_));
 sky130_fd_sc_hd__nand2_1 _23974_ (.A(_04153_),
    .B(_04154_),
    .Y(_04155_));
 sky130_fd_sc_hd__buf_2 _23975_ (.A(_03764_),
    .X(_04156_));
 sky130_fd_sc_hd__nand2_1 _23976_ (.A(_04156_),
    .B(_04052_),
    .Y(_04157_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _23977_ (.A(_02567_),
    .X(_04158_));
 sky130_fd_sc_hd__a21oi_1 _23978_ (.A1(_04157_),
    .A2(_04054_),
    .B1(_04158_),
    .Y(_04159_));
 sky130_fd_sc_hd__and3_1 _23979_ (.A(_02567_),
    .B(_04157_),
    .C(_04054_),
    .X(_04160_));
 sky130_fd_sc_hd__or2_1 _23980_ (.A(_04159_),
    .B(_04160_),
    .X(_04161_));
 sky130_fd_sc_hd__xor2_1 _23981_ (.A(_04155_),
    .B(_04161_),
    .X(_04162_));
 sky130_fd_sc_hd__o21ba_1 _23982_ (.A1(_04057_),
    .A2(_04059_),
    .B1_N(_04066_),
    .X(_04163_));
 sky130_fd_sc_hd__xnor2_1 _23983_ (.A(_04162_),
    .B(_04163_),
    .Y(_04164_));
 sky130_fd_sc_hd__nand2_1 _23984_ (.A(_04063_),
    .B(_04164_),
    .Y(_04165_));
 sky130_fd_sc_hd__or2_1 _23985_ (.A(_04063_),
    .B(_04164_),
    .X(_04166_));
 sky130_fd_sc_hd__nand2_1 _23986_ (.A(_04165_),
    .B(_04166_),
    .Y(_04167_));
 sky130_fd_sc_hd__a21oi_1 _23987_ (.A1(_04078_),
    .A2(_04071_),
    .B1(_04167_),
    .Y(_04168_));
 sky130_fd_sc_hd__and3_1 _23988_ (.A(_04078_),
    .B(_04071_),
    .C(_04167_),
    .X(_04169_));
 sky130_fd_sc_hd__nor2_2 _23989_ (.A(_04168_),
    .B(_04169_),
    .Y(_04170_));
 sky130_fd_sc_hd__or2_1 _23990_ (.A(_03977_),
    .B(_04074_),
    .X(_04171_));
 sky130_fd_sc_hd__and3_1 _23991_ (.A(_03983_),
    .B(_04075_),
    .C(_04171_),
    .X(_04172_));
 sky130_fd_sc_hd__a21o_1 _23992_ (.A1(_03978_),
    .A2(_04075_),
    .B1(_04074_),
    .X(_04173_));
 sky130_fd_sc_hd__a21oi_4 _23993_ (.A1(_03982_),
    .A2(_04172_),
    .B1(_04173_),
    .Y(_04174_));
 sky130_fd_sc_hd__xor2_4 _23994_ (.A(_04170_),
    .B(_04174_),
    .X(_00102_));
 sky130_fd_sc_hd__or2b_1 _23995_ (.A(_04163_),
    .B_N(_04162_),
    .X(_04175_));
 sky130_fd_sc_hd__and2b_1 _23996_ (.A_N(_14262_),
    .B(_13804_),
    .X(_04176_));
 sky130_fd_sc_hd__a21oi_1 _23997_ (.A1(_02472_),
    .A2(_04079_),
    .B1(_04176_),
    .Y(_04177_));
 sky130_fd_sc_hd__and3_1 _23998_ (.A(_13869_),
    .B(_04079_),
    .C(_04176_),
    .X(_04178_));
 sky130_fd_sc_hd__nor2_1 _23999_ (.A(_04177_),
    .B(_04178_),
    .Y(_04179_));
 sky130_fd_sc_hd__nand2_1 _24000_ (.A(_04092_),
    .B(_04084_),
    .Y(_04180_));
 sky130_fd_sc_hd__xnor2_1 _24001_ (.A(_04179_),
    .B(_04180_),
    .Y(_04181_));
 sky130_fd_sc_hd__o21ba_1 _24002_ (.A1(_04081_),
    .A2(_04085_),
    .B1_N(_04082_),
    .X(_04182_));
 sky130_fd_sc_hd__xnor2_1 _24003_ (.A(_04181_),
    .B(_04182_),
    .Y(_04183_));
 sky130_fd_sc_hd__a22oi_1 _24004_ (.A1(_04090_),
    .A2(_04095_),
    .B1(_13816_),
    .B2(_04094_),
    .Y(_04184_));
 sky130_fd_sc_hd__and4_1 _24005_ (.A(_04094_),
    .B(_01718_),
    .C(_04095_),
    .D(_13815_),
    .X(_04185_));
 sky130_fd_sc_hd__or2_1 _24006_ (.A(_04184_),
    .B(_04185_),
    .X(_04186_));
 sky130_fd_sc_hd__nand2_1 _24007_ (.A(_03804_),
    .B(_13819_),
    .Y(_04187_));
 sky130_fd_sc_hd__xor2_1 _24008_ (.A(_04186_),
    .B(_04187_),
    .X(_04188_));
 sky130_fd_sc_hd__xnor2_1 _24009_ (.A(_04183_),
    .B(_04188_),
    .Y(_04189_));
 sky130_fd_sc_hd__and2b_1 _24010_ (.A_N(_04087_),
    .B(_04086_),
    .X(_04190_));
 sky130_fd_sc_hd__a21oi_1 _24011_ (.A1(_04088_),
    .A2(_04100_),
    .B1(_04190_),
    .Y(_04191_));
 sky130_fd_sc_hd__xor2_1 _24012_ (.A(_04189_),
    .B(_04191_),
    .X(_04192_));
 sky130_fd_sc_hd__o21ba_1 _24013_ (.A1(_04106_),
    .A2(_04109_),
    .B1_N(_04107_),
    .X(_04193_));
 sky130_fd_sc_hd__o21ba_1 _24014_ (.A1(_04093_),
    .A2(_04099_),
    .B1_N(_04096_),
    .X(_04194_));
 sky130_fd_sc_hd__a22o_1 _24015_ (.A1(_03609_),
    .A2(_03628_),
    .B1(_14564_),
    .B2(_12773_),
    .X(_04195_));
 sky130_fd_sc_hd__and3_1 _24016_ (.A(_12773_),
    .B(_03609_),
    .C(_14038_),
    .X(_04196_));
 sky130_fd_sc_hd__nand2_1 _24017_ (.A(_03628_),
    .B(_04196_),
    .Y(_04197_));
 sky130_fd_sc_hd__nand2_1 _24018_ (.A(_04195_),
    .B(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__xor2_1 _24019_ (.A(_04109_),
    .B(_04198_),
    .X(_04199_));
 sky130_fd_sc_hd__xnor2_1 _24020_ (.A(_04194_),
    .B(_04199_),
    .Y(_04200_));
 sky130_fd_sc_hd__xnor2_1 _24021_ (.A(_04193_),
    .B(_04200_),
    .Y(_04201_));
 sky130_fd_sc_hd__xnor2_1 _24022_ (.A(_04192_),
    .B(_04201_),
    .Y(_04202_));
 sky130_fd_sc_hd__nor2_1 _24023_ (.A(_04101_),
    .B(_04103_),
    .Y(_04203_));
 sky130_fd_sc_hd__a21oi_1 _24024_ (.A1(_04104_),
    .A2(_04116_),
    .B1(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__xnor2_1 _24025_ (.A(_04202_),
    .B(_04204_),
    .Y(_04205_));
 sky130_fd_sc_hd__a21oi_1 _24026_ (.A1(_03826_),
    .A2(_04122_),
    .B1(_04120_),
    .Y(_04206_));
 sky130_fd_sc_hd__a21o_1 _24027_ (.A1(_04111_),
    .A2(_04114_),
    .B1(_04124_),
    .X(_04207_));
 sky130_fd_sc_hd__clkbuf_2 _24028_ (.A(_04124_),
    .X(_04208_));
 sky130_fd_sc_hd__nand3_1 _24029_ (.A(_04111_),
    .B(_04114_),
    .C(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__nand2_1 _24030_ (.A(_04207_),
    .B(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hd__xnor2_1 _24031_ (.A(_04206_),
    .B(_04210_),
    .Y(_04211_));
 sky130_fd_sc_hd__nor2_1 _24032_ (.A(_04205_),
    .B(_04211_),
    .Y(_04212_));
 sky130_fd_sc_hd__and2_1 _24033_ (.A(_04205_),
    .B(_04211_),
    .X(_04213_));
 sky130_fd_sc_hd__or2_1 _24034_ (.A(_04212_),
    .B(_04213_),
    .X(_04214_));
 sky130_fd_sc_hd__nor2_1 _24035_ (.A(_04117_),
    .B(_04118_),
    .Y(_04215_));
 sky130_fd_sc_hd__a21oi_1 _24036_ (.A1(_04119_),
    .A2(_04128_),
    .B1(_04215_),
    .Y(_04216_));
 sky130_fd_sc_hd__xor2_1 _24037_ (.A(_04214_),
    .B(_04216_),
    .X(_04217_));
 sky130_fd_sc_hd__and2b_1 _24038_ (.A_N(_04121_),
    .B(_04127_),
    .X(_04218_));
 sky130_fd_sc_hd__nor2_1 _24039_ (.A(_04125_),
    .B(_04218_),
    .Y(_04219_));
 sky130_fd_sc_hd__xnor2_1 _24040_ (.A(_04044_),
    .B(_04219_),
    .Y(_04220_));
 sky130_fd_sc_hd__or2_1 _24041_ (.A(_04040_),
    .B(_04220_),
    .X(_04221_));
 sky130_fd_sc_hd__clkbuf_2 _24042_ (.A(_04040_),
    .X(_04222_));
 sky130_fd_sc_hd__nand2_1 _24043_ (.A(_04222_),
    .B(_04220_),
    .Y(_04223_));
 sky130_fd_sc_hd__and2_1 _24044_ (.A(_04221_),
    .B(_04223_),
    .X(_04224_));
 sky130_fd_sc_hd__xnor2_1 _24045_ (.A(_04217_),
    .B(_04224_),
    .Y(_04225_));
 sky130_fd_sc_hd__nor2_1 _24046_ (.A(_04129_),
    .B(_04132_),
    .Y(_04226_));
 sky130_fd_sc_hd__a21oi_1 _24047_ (.A1(_04133_),
    .A2(_04139_),
    .B1(_04226_),
    .Y(_04227_));
 sky130_fd_sc_hd__xor2_1 _24048_ (.A(_04225_),
    .B(_04227_),
    .X(_04228_));
 sky130_fd_sc_hd__clkbuf_2 _24049_ (.A(_04044_),
    .X(_04229_));
 sky130_fd_sc_hd__o21a_1 _24050_ (.A1(_04229_),
    .A2(_04135_),
    .B1(_04137_),
    .X(_04230_));
 sky130_fd_sc_hd__xnor2_1 _24051_ (.A(_03764_),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__nand2_1 _24052_ (.A(_03773_),
    .B(_04231_),
    .Y(_04232_));
 sky130_fd_sc_hd__or2_1 _24053_ (.A(_03773_),
    .B(_04231_),
    .X(_04233_));
 sky130_fd_sc_hd__and2_1 _24054_ (.A(_04232_),
    .B(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__xnor2_1 _24055_ (.A(_04228_),
    .B(_04234_),
    .Y(_04235_));
 sky130_fd_sc_hd__nor2_1 _24056_ (.A(_04140_),
    .B(_04143_),
    .Y(_04236_));
 sky130_fd_sc_hd__a21oi_1 _24057_ (.A1(_04144_),
    .A2(_04149_),
    .B1(_04236_),
    .Y(_04237_));
 sky130_fd_sc_hd__xnor2_1 _24058_ (.A(_04235_),
    .B(_04237_),
    .Y(_04238_));
 sky130_fd_sc_hd__or3_1 _24059_ (.A(_03471_),
    .B(_03472_),
    .C(_04145_),
    .X(_04239_));
 sky130_fd_sc_hd__a21oi_1 _24060_ (.A1(_04239_),
    .A2(_04147_),
    .B1(_02567_),
    .Y(_04240_));
 sky130_fd_sc_hd__and3_1 _24061_ (.A(_02567_),
    .B(_04239_),
    .C(_04147_),
    .X(_04241_));
 sky130_fd_sc_hd__or2_1 _24062_ (.A(_04240_),
    .B(_04241_),
    .X(_04242_));
 sky130_fd_sc_hd__xor2_1 _24063_ (.A(_04238_),
    .B(_04242_),
    .X(_04243_));
 sky130_fd_sc_hd__o21a_1 _24064_ (.A1(_04155_),
    .A2(_04161_),
    .B1(_04153_),
    .X(_04244_));
 sky130_fd_sc_hd__xnor2_1 _24065_ (.A(_04243_),
    .B(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__nand2_1 _24066_ (.A(_04159_),
    .B(_04245_),
    .Y(_04246_));
 sky130_fd_sc_hd__or2_1 _24067_ (.A(_04159_),
    .B(_04245_),
    .X(_04247_));
 sky130_fd_sc_hd__nand2_1 _24068_ (.A(_04246_),
    .B(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__and3_1 _24069_ (.A(_04175_),
    .B(_04165_),
    .C(_04248_),
    .X(_04249_));
 sky130_fd_sc_hd__a21oi_1 _24070_ (.A1(_04175_),
    .A2(_04165_),
    .B1(_04248_),
    .Y(_04250_));
 sky130_fd_sc_hd__nor2_1 _24071_ (.A(_04249_),
    .B(_04250_),
    .Y(_04251_));
 sky130_fd_sc_hd__a21oi_1 _24072_ (.A1(_04170_),
    .A2(_04174_),
    .B1(_04168_),
    .Y(_04252_));
 sky130_fd_sc_hd__xnor2_1 _24073_ (.A(_04251_),
    .B(_04252_),
    .Y(_00103_));
 sky130_fd_sc_hd__or2b_1 _24074_ (.A(_04244_),
    .B_N(_04243_),
    .X(_04253_));
 sky130_fd_sc_hd__buf_2 _24075_ (.A(_04079_),
    .X(_04254_));
 sky130_fd_sc_hd__and2b_1 _24076_ (.A_N(_13869_),
    .B(_13805_),
    .X(_04255_));
 sky130_fd_sc_hd__a21oi_1 _24077_ (.A1(_04092_),
    .A2(_04254_),
    .B1(_04255_),
    .Y(_04256_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _24078_ (.A(_04079_),
    .X(_04257_));
 sky130_fd_sc_hd__and3_1 _24079_ (.A(_04092_),
    .B(_04257_),
    .C(_04255_),
    .X(_04258_));
 sky130_fd_sc_hd__nor2_1 _24080_ (.A(_04256_),
    .B(_04258_),
    .Y(_04259_));
 sky130_fd_sc_hd__nand2_1 _24081_ (.A(_04090_),
    .B(_04084_),
    .Y(_04260_));
 sky130_fd_sc_hd__xnor2_2 _24082_ (.A(_04259_),
    .B(_04260_),
    .Y(_04261_));
 sky130_fd_sc_hd__o21ba_1 _24083_ (.A1(_04177_),
    .A2(_04180_),
    .B1_N(_04178_),
    .X(_04262_));
 sky130_fd_sc_hd__xnor2_2 _24084_ (.A(_04261_),
    .B(_04262_),
    .Y(_04263_));
 sky130_fd_sc_hd__clkbuf_2 _24085_ (.A(_13825_),
    .X(_04264_));
 sky130_fd_sc_hd__a22oi_1 _24086_ (.A1(_04095_),
    .A2(_04264_),
    .B1(_13818_),
    .B2(_04089_),
    .Y(_04265_));
 sky130_fd_sc_hd__and4_1 _24087_ (.A(_04094_),
    .B(_04095_),
    .C(_04264_),
    .D(_13818_),
    .X(_04266_));
 sky130_fd_sc_hd__nor2_1 _24088_ (.A(_04265_),
    .B(_04266_),
    .Y(_04267_));
 sky130_fd_sc_hd__nand2_1 _24089_ (.A(_04098_),
    .B(_14214_),
    .Y(_04268_));
 sky130_fd_sc_hd__xnor2_2 _24090_ (.A(_04267_),
    .B(_04268_),
    .Y(_04269_));
 sky130_fd_sc_hd__xnor2_2 _24091_ (.A(_04263_),
    .B(_04269_),
    .Y(_04270_));
 sky130_fd_sc_hd__and2b_1 _24092_ (.A_N(_04182_),
    .B(_04181_),
    .X(_04271_));
 sky130_fd_sc_hd__a21oi_1 _24093_ (.A1(_04183_),
    .A2(_04188_),
    .B1(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__xor2_1 _24094_ (.A(_04270_),
    .B(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__o21ai_1 _24095_ (.A1(_04109_),
    .A2(_04198_),
    .B1(_04197_),
    .Y(_04274_));
 sky130_fd_sc_hd__nor2_1 _24096_ (.A(_04186_),
    .B(_04187_),
    .Y(_04275_));
 sky130_fd_sc_hd__o21ai_1 _24097_ (.A1(_12773_),
    .A2(_03609_),
    .B1(_14563_),
    .Y(_04276_));
 sky130_fd_sc_hd__nor2_1 _24098_ (.A(_04196_),
    .B(_04276_),
    .Y(_04277_));
 sky130_fd_sc_hd__xnor2_2 _24099_ (.A(_04109_),
    .B(_04277_),
    .Y(_04278_));
 sky130_fd_sc_hd__o21a_1 _24100_ (.A1(_04185_),
    .A2(_04275_),
    .B1(_04278_),
    .X(_04279_));
 sky130_fd_sc_hd__nor3_1 _24101_ (.A(_04185_),
    .B(_04275_),
    .C(_04278_),
    .Y(_04280_));
 sky130_fd_sc_hd__nor2_1 _24102_ (.A(_04279_),
    .B(_04280_),
    .Y(_04281_));
 sky130_fd_sc_hd__xor2_1 _24103_ (.A(_04274_),
    .B(_04281_),
    .X(_04282_));
 sky130_fd_sc_hd__xnor2_1 _24104_ (.A(_04273_),
    .B(_04282_),
    .Y(_04283_));
 sky130_fd_sc_hd__nor2_1 _24105_ (.A(_04189_),
    .B(_04191_),
    .Y(_04284_));
 sky130_fd_sc_hd__a21oi_1 _24106_ (.A1(_04192_),
    .A2(_04201_),
    .B1(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__xnor2_1 _24107_ (.A(_04283_),
    .B(_04285_),
    .Y(_04286_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _24108_ (.A(_04206_),
    .X(_04287_));
 sky130_fd_sc_hd__and2b_1 _24109_ (.A_N(_04194_),
    .B(_04199_),
    .X(_04288_));
 sky130_fd_sc_hd__and2b_1 _24110_ (.A_N(_04193_),
    .B(_04200_),
    .X(_04289_));
 sky130_fd_sc_hd__nor2_1 _24111_ (.A(_04288_),
    .B(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__xnor2_1 _24112_ (.A(_04208_),
    .B(_04290_),
    .Y(_04291_));
 sky130_fd_sc_hd__xnor2_1 _24113_ (.A(_04287_),
    .B(_04291_),
    .Y(_04292_));
 sky130_fd_sc_hd__nor2_1 _24114_ (.A(_04286_),
    .B(_04292_),
    .Y(_04293_));
 sky130_fd_sc_hd__and2_1 _24115_ (.A(_04286_),
    .B(_04292_),
    .X(_04294_));
 sky130_fd_sc_hd__nor2_1 _24116_ (.A(_04293_),
    .B(_04294_),
    .Y(_04295_));
 sky130_fd_sc_hd__o21ba_1 _24117_ (.A1(_04202_),
    .A2(_04204_),
    .B1_N(_04212_),
    .X(_04296_));
 sky130_fd_sc_hd__xnor2_1 _24118_ (.A(_04295_),
    .B(_04296_),
    .Y(_04297_));
 sky130_fd_sc_hd__clkbuf_2 _24119_ (.A(_04040_),
    .X(_04298_));
 sky130_fd_sc_hd__clkbuf_2 _24120_ (.A(_04287_),
    .X(_04299_));
 sky130_fd_sc_hd__o21a_1 _24121_ (.A1(_04299_),
    .A2(_04210_),
    .B1(_04207_),
    .X(_04300_));
 sky130_fd_sc_hd__or2_1 _24122_ (.A(_04229_),
    .B(_04300_),
    .X(_04301_));
 sky130_fd_sc_hd__nand2_1 _24123_ (.A(_04229_),
    .B(_04300_),
    .Y(_04302_));
 sky130_fd_sc_hd__nand2_1 _24124_ (.A(_04301_),
    .B(_04302_),
    .Y(_04303_));
 sky130_fd_sc_hd__xor2_1 _24125_ (.A(_04298_),
    .B(_04303_),
    .X(_04304_));
 sky130_fd_sc_hd__nand2_1 _24126_ (.A(_04297_),
    .B(_04304_),
    .Y(_04305_));
 sky130_fd_sc_hd__or2_1 _24127_ (.A(_04297_),
    .B(_04304_),
    .X(_04306_));
 sky130_fd_sc_hd__nand2_1 _24128_ (.A(_04305_),
    .B(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__nor2_1 _24129_ (.A(_04214_),
    .B(_04216_),
    .Y(_04308_));
 sky130_fd_sc_hd__a21oi_1 _24130_ (.A1(_04217_),
    .A2(_04224_),
    .B1(_04308_),
    .Y(_04309_));
 sky130_fd_sc_hd__xor2_1 _24131_ (.A(_04307_),
    .B(_04309_),
    .X(_04310_));
 sky130_fd_sc_hd__clkbuf_2 _24132_ (.A(_03874_),
    .X(_04311_));
 sky130_fd_sc_hd__clkbuf_2 _24133_ (.A(_04229_),
    .X(_04312_));
 sky130_fd_sc_hd__o21a_1 _24134_ (.A1(_04312_),
    .A2(_04219_),
    .B1(_04221_),
    .X(_04313_));
 sky130_fd_sc_hd__xnor2_1 _24135_ (.A(_04156_),
    .B(_04313_),
    .Y(_04314_));
 sky130_fd_sc_hd__nand2_1 _24136_ (.A(_04311_),
    .B(_04314_),
    .Y(_04315_));
 sky130_fd_sc_hd__or2_1 _24137_ (.A(_03874_),
    .B(_04314_),
    .X(_04316_));
 sky130_fd_sc_hd__and2_1 _24138_ (.A(_04315_),
    .B(_04316_),
    .X(_04317_));
 sky130_fd_sc_hd__xnor2_1 _24139_ (.A(_04310_),
    .B(_04317_),
    .Y(_04318_));
 sky130_fd_sc_hd__nor2_1 _24140_ (.A(_04225_),
    .B(_04227_),
    .Y(_04319_));
 sky130_fd_sc_hd__a21oi_1 _24141_ (.A1(_04228_),
    .A2(_04234_),
    .B1(_04319_),
    .Y(_04320_));
 sky130_fd_sc_hd__xnor2_1 _24142_ (.A(_04318_),
    .B(_04320_),
    .Y(_04321_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _24143_ (.A(_03471_),
    .X(_04322_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _24144_ (.A(_03472_),
    .X(_04323_));
 sky130_fd_sc_hd__or3_1 _24145_ (.A(_04322_),
    .B(_04323_),
    .C(_04230_),
    .X(_04324_));
 sky130_fd_sc_hd__a21oi_1 _24146_ (.A1(_04324_),
    .A2(_04232_),
    .B1(_04158_),
    .Y(_04325_));
 sky130_fd_sc_hd__and3_1 _24147_ (.A(_04158_),
    .B(_04324_),
    .C(_04232_),
    .X(_04326_));
 sky130_fd_sc_hd__or2_1 _24148_ (.A(_04325_),
    .B(_04326_),
    .X(_04327_));
 sky130_fd_sc_hd__xor2_1 _24149_ (.A(_04321_),
    .B(_04327_),
    .X(_04328_));
 sky130_fd_sc_hd__or2_1 _24150_ (.A(_04235_),
    .B(_04237_),
    .X(_04329_));
 sky130_fd_sc_hd__o21a_1 _24151_ (.A1(_04238_),
    .A2(_04242_),
    .B1(_04329_),
    .X(_04330_));
 sky130_fd_sc_hd__xnor2_1 _24152_ (.A(_04328_),
    .B(_04330_),
    .Y(_04331_));
 sky130_fd_sc_hd__nand2_1 _24153_ (.A(_04240_),
    .B(_04331_),
    .Y(_04332_));
 sky130_fd_sc_hd__or2_1 _24154_ (.A(_04240_),
    .B(_04331_),
    .X(_04333_));
 sky130_fd_sc_hd__nand2_1 _24155_ (.A(_04332_),
    .B(_04333_),
    .Y(_04334_));
 sky130_fd_sc_hd__a21oi_1 _24156_ (.A1(_04253_),
    .A2(_04246_),
    .B1(_04334_),
    .Y(_04335_));
 sky130_fd_sc_hd__nand3_1 _24157_ (.A(_04253_),
    .B(_04246_),
    .C(_04334_),
    .Y(_04336_));
 sky130_fd_sc_hd__or2b_1 _24158_ (.A(_04335_),
    .B_N(_04336_),
    .X(_04337_));
 sky130_fd_sc_hd__nor2_1 _24159_ (.A(_04168_),
    .B(_04250_),
    .Y(_04338_));
 sky130_fd_sc_hd__nor2_1 _24160_ (.A(_04249_),
    .B(_04338_),
    .Y(_04339_));
 sky130_fd_sc_hd__a31o_1 _24161_ (.A1(_04170_),
    .A2(_04174_),
    .A3(_04251_),
    .B1(_04339_),
    .X(_04340_));
 sky130_fd_sc_hd__xnor2_1 _24162_ (.A(_04337_),
    .B(_04340_),
    .Y(_00104_));
 sky130_fd_sc_hd__or2b_1 _24163_ (.A(_04330_),
    .B_N(_04328_),
    .X(_04341_));
 sky130_fd_sc_hd__and2b_1 _24164_ (.A_N(_02610_),
    .B(_13804_),
    .X(_04342_));
 sky130_fd_sc_hd__a21oi_1 _24165_ (.A1(_04090_),
    .A2(_04257_),
    .B1(_04342_),
    .Y(_04343_));
 sky130_fd_sc_hd__and3_1 _24166_ (.A(_01718_),
    .B(_04257_),
    .C(_04342_),
    .X(_04344_));
 sky130_fd_sc_hd__nor2_1 _24167_ (.A(_04343_),
    .B(_04344_),
    .Y(_04345_));
 sky130_fd_sc_hd__nand2_1 _24168_ (.A(_13816_),
    .B(_04084_),
    .Y(_04346_));
 sky130_fd_sc_hd__xnor2_1 _24169_ (.A(_04345_),
    .B(_04346_),
    .Y(_04347_));
 sky130_fd_sc_hd__o21ba_1 _24170_ (.A1(_04256_),
    .A2(_04260_),
    .B1_N(_04258_),
    .X(_04348_));
 sky130_fd_sc_hd__xor2_1 _24171_ (.A(_04347_),
    .B(_04348_),
    .X(_04349_));
 sky130_fd_sc_hd__a22oi_1 _24172_ (.A1(_04091_),
    .A2(_13818_),
    .B1(_03628_),
    .B2(_04089_),
    .Y(_04350_));
 sky130_fd_sc_hd__and4_1 _24173_ (.A(_04089_),
    .B(_04091_),
    .C(_13818_),
    .D(_03628_),
    .X(_04351_));
 sky130_fd_sc_hd__nor2_1 _24174_ (.A(_04350_),
    .B(_04351_),
    .Y(_04352_));
 sky130_fd_sc_hd__nand2_2 _24175_ (.A(_03804_),
    .B(_14564_),
    .Y(_04353_));
 sky130_fd_sc_hd__xor2_1 _24176_ (.A(_04352_),
    .B(_04353_),
    .X(_04354_));
 sky130_fd_sc_hd__xnor2_1 _24177_ (.A(_04349_),
    .B(_04354_),
    .Y(_04355_));
 sky130_fd_sc_hd__and2b_1 _24178_ (.A_N(_04262_),
    .B(_04261_),
    .X(_04356_));
 sky130_fd_sc_hd__a21oi_2 _24179_ (.A1(_04263_),
    .A2(_04269_),
    .B1(_04356_),
    .Y(_04357_));
 sky130_fd_sc_hd__xnor2_1 _24180_ (.A(_04355_),
    .B(_04357_),
    .Y(_04358_));
 sky130_fd_sc_hd__o21bai_1 _24181_ (.A1(_04109_),
    .A2(_04276_),
    .B1_N(_04196_),
    .Y(_04359_));
 sky130_fd_sc_hd__a31o_1 _24182_ (.A1(_04098_),
    .A2(_14213_),
    .A3(_04267_),
    .B1(_04266_),
    .X(_04360_));
 sky130_fd_sc_hd__xor2_1 _24183_ (.A(_04278_),
    .B(_04360_),
    .X(_04361_));
 sky130_fd_sc_hd__and2_1 _24184_ (.A(_04359_),
    .B(_04361_),
    .X(_04362_));
 sky130_fd_sc_hd__clkbuf_2 _24185_ (.A(_04359_),
    .X(_04363_));
 sky130_fd_sc_hd__nor2_1 _24186_ (.A(_04363_),
    .B(_04361_),
    .Y(_04364_));
 sky130_fd_sc_hd__or2_1 _24187_ (.A(_04362_),
    .B(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__xnor2_1 _24188_ (.A(_04358_),
    .B(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hd__nor2_1 _24189_ (.A(_04270_),
    .B(_04272_),
    .Y(_04367_));
 sky130_fd_sc_hd__a21oi_1 _24190_ (.A1(_04273_),
    .A2(_04282_),
    .B1(_04367_),
    .Y(_04368_));
 sky130_fd_sc_hd__xnor2_1 _24191_ (.A(_04366_),
    .B(_04368_),
    .Y(_04369_));
 sky130_fd_sc_hd__a21oi_1 _24192_ (.A1(_04274_),
    .A2(_04281_),
    .B1(_04279_),
    .Y(_04370_));
 sky130_fd_sc_hd__xnor2_1 _24193_ (.A(_04124_),
    .B(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hd__or2_1 _24194_ (.A(_04206_),
    .B(_04371_),
    .X(_04372_));
 sky130_fd_sc_hd__nand2_1 _24195_ (.A(_04287_),
    .B(_04371_),
    .Y(_04373_));
 sky130_fd_sc_hd__nand2_1 _24196_ (.A(_04372_),
    .B(_04373_),
    .Y(_04374_));
 sky130_fd_sc_hd__nor2_1 _24197_ (.A(_04369_),
    .B(_04374_),
    .Y(_04375_));
 sky130_fd_sc_hd__and2_1 _24198_ (.A(_04369_),
    .B(_04374_),
    .X(_04376_));
 sky130_fd_sc_hd__nor2_1 _24199_ (.A(_04375_),
    .B(_04376_),
    .Y(_04377_));
 sky130_fd_sc_hd__o21ba_1 _24200_ (.A1(_04283_),
    .A2(_04285_),
    .B1_N(_04293_),
    .X(_04378_));
 sky130_fd_sc_hd__xnor2_1 _24201_ (.A(_04377_),
    .B(_04378_),
    .Y(_04379_));
 sky130_fd_sc_hd__or2_1 _24202_ (.A(_04208_),
    .B(_04290_),
    .X(_04380_));
 sky130_fd_sc_hd__o21a_1 _24203_ (.A1(_04287_),
    .A2(_04291_),
    .B1(_04380_),
    .X(_04381_));
 sky130_fd_sc_hd__or2_1 _24204_ (.A(_04044_),
    .B(_04381_),
    .X(_04382_));
 sky130_fd_sc_hd__nand2_1 _24205_ (.A(_04229_),
    .B(_04381_),
    .Y(_04383_));
 sky130_fd_sc_hd__nand2_1 _24206_ (.A(_04382_),
    .B(_04383_),
    .Y(_04384_));
 sky130_fd_sc_hd__xor2_1 _24207_ (.A(_04222_),
    .B(_04384_),
    .X(_04385_));
 sky130_fd_sc_hd__nand2_1 _24208_ (.A(_04379_),
    .B(_04385_),
    .Y(_04386_));
 sky130_fd_sc_hd__or2_1 _24209_ (.A(_04379_),
    .B(_04385_),
    .X(_04387_));
 sky130_fd_sc_hd__nand2_1 _24210_ (.A(_04386_),
    .B(_04387_),
    .Y(_04388_));
 sky130_fd_sc_hd__o31a_1 _24211_ (.A1(_04293_),
    .A2(_04294_),
    .A3(_04296_),
    .B1(_04305_),
    .X(_04389_));
 sky130_fd_sc_hd__nor2_1 _24212_ (.A(_04388_),
    .B(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__and2_1 _24213_ (.A(_04388_),
    .B(_04389_),
    .X(_04391_));
 sky130_fd_sc_hd__nor2_1 _24214_ (.A(_04390_),
    .B(_04391_),
    .Y(_04392_));
 sky130_fd_sc_hd__o21a_1 _24215_ (.A1(_04298_),
    .A2(_04303_),
    .B1(_04301_),
    .X(_04393_));
 sky130_fd_sc_hd__xnor2_1 _24216_ (.A(_04156_),
    .B(_04393_),
    .Y(_04394_));
 sky130_fd_sc_hd__nand2_1 _24217_ (.A(_04311_),
    .B(_04394_),
    .Y(_04395_));
 sky130_fd_sc_hd__or2_1 _24218_ (.A(_03874_),
    .B(_04394_),
    .X(_04396_));
 sky130_fd_sc_hd__and2_1 _24219_ (.A(_04395_),
    .B(_04396_),
    .X(_04397_));
 sky130_fd_sc_hd__xnor2_1 _24220_ (.A(_04392_),
    .B(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__nor2_1 _24221_ (.A(_04307_),
    .B(_04309_),
    .Y(_04399_));
 sky130_fd_sc_hd__a21oi_1 _24222_ (.A1(_04310_),
    .A2(_04317_),
    .B1(_04399_),
    .Y(_04400_));
 sky130_fd_sc_hd__xnor2_1 _24223_ (.A(_04398_),
    .B(_04400_),
    .Y(_04401_));
 sky130_fd_sc_hd__or3_1 _24224_ (.A(_04322_),
    .B(_04323_),
    .C(_04313_),
    .X(_04402_));
 sky130_fd_sc_hd__a21oi_1 _24225_ (.A1(_04402_),
    .A2(_04315_),
    .B1(_04158_),
    .Y(_04403_));
 sky130_fd_sc_hd__and3_1 _24226_ (.A(_04158_),
    .B(_04402_),
    .C(_04315_),
    .X(_04404_));
 sky130_fd_sc_hd__or2_1 _24227_ (.A(_04403_),
    .B(_04404_),
    .X(_04405_));
 sky130_fd_sc_hd__nor2_1 _24228_ (.A(_04401_),
    .B(_04405_),
    .Y(_04406_));
 sky130_fd_sc_hd__and2_1 _24229_ (.A(_04401_),
    .B(_04405_),
    .X(_04407_));
 sky130_fd_sc_hd__nor2_1 _24230_ (.A(_04406_),
    .B(_04407_),
    .Y(_04408_));
 sky130_fd_sc_hd__or2_1 _24231_ (.A(_04318_),
    .B(_04320_),
    .X(_04409_));
 sky130_fd_sc_hd__o21a_1 _24232_ (.A1(_04321_),
    .A2(_04327_),
    .B1(_04409_),
    .X(_04410_));
 sky130_fd_sc_hd__xnor2_1 _24233_ (.A(_04408_),
    .B(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hd__xnor2_1 _24234_ (.A(_04325_),
    .B(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__nand3_1 _24235_ (.A(_04341_),
    .B(_04332_),
    .C(_04412_),
    .Y(_04413_));
 sky130_vsdinv _24236_ (.A(_04413_),
    .Y(_04414_));
 sky130_fd_sc_hd__a21oi_1 _24237_ (.A1(_04341_),
    .A2(_04332_),
    .B1(_04412_),
    .Y(_04415_));
 sky130_fd_sc_hd__nor2_1 _24238_ (.A(_04414_),
    .B(_04415_),
    .Y(_04416_));
 sky130_fd_sc_hd__a21oi_1 _24239_ (.A1(_04336_),
    .A2(_04340_),
    .B1(_04335_),
    .Y(_04417_));
 sky130_fd_sc_hd__xnor2_1 _24240_ (.A(_04416_),
    .B(_04417_),
    .Y(_00105_));
 sky130_fd_sc_hd__or3_1 _24241_ (.A(_04406_),
    .B(_04407_),
    .C(_04410_),
    .X(_04418_));
 sky130_fd_sc_hd__nand2_1 _24242_ (.A(_04325_),
    .B(_04411_),
    .Y(_04419_));
 sky130_fd_sc_hd__and2b_1 _24243_ (.A_N(_01844_),
    .B(_13804_),
    .X(_04420_));
 sky130_fd_sc_hd__a21oi_1 _24244_ (.A1(_04264_),
    .A2(_04254_),
    .B1(_04420_),
    .Y(_04421_));
 sky130_fd_sc_hd__and3_1 _24245_ (.A(_04264_),
    .B(_04257_),
    .C(_04420_),
    .X(_04422_));
 sky130_fd_sc_hd__nor2_1 _24246_ (.A(_04421_),
    .B(_04422_),
    .Y(_04423_));
 sky130_fd_sc_hd__nand2_1 _24247_ (.A(_04084_),
    .B(_13819_),
    .Y(_04424_));
 sky130_fd_sc_hd__xnor2_1 _24248_ (.A(_04423_),
    .B(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hd__o21ba_1 _24249_ (.A1(_04343_),
    .A2(_04346_),
    .B1_N(_04344_),
    .X(_04426_));
 sky130_fd_sc_hd__xor2_1 _24250_ (.A(_04425_),
    .B(_04426_),
    .X(_04427_));
 sky130_fd_sc_hd__a22oi_2 _24251_ (.A1(_04091_),
    .A2(_14213_),
    .B1(_14564_),
    .B2(_04089_),
    .Y(_04428_));
 sky130_fd_sc_hd__and3_1 _24252_ (.A(_04094_),
    .B(_04095_),
    .C(_14563_),
    .X(_04429_));
 sky130_fd_sc_hd__and2_1 _24253_ (.A(_14213_),
    .B(_04429_),
    .X(_04430_));
 sky130_fd_sc_hd__nor3_1 _24254_ (.A(_04353_),
    .B(_04428_),
    .C(_04430_),
    .Y(_04431_));
 sky130_fd_sc_hd__o21a_1 _24255_ (.A1(_04428_),
    .A2(_04430_),
    .B1(_04353_),
    .X(_04432_));
 sky130_fd_sc_hd__nor2_1 _24256_ (.A(_04431_),
    .B(_04432_),
    .Y(_04433_));
 sky130_fd_sc_hd__xnor2_1 _24257_ (.A(_04427_),
    .B(_04433_),
    .Y(_04434_));
 sky130_fd_sc_hd__or2b_1 _24258_ (.A(_04348_),
    .B_N(_04347_),
    .X(_04435_));
 sky130_fd_sc_hd__o21a_1 _24259_ (.A1(_04349_),
    .A2(_04354_),
    .B1(_04435_),
    .X(_04436_));
 sky130_fd_sc_hd__xor2_1 _24260_ (.A(_04434_),
    .B(_04436_),
    .X(_04437_));
 sky130_fd_sc_hd__a31o_1 _24261_ (.A1(_04098_),
    .A2(_14565_),
    .A3(_04352_),
    .B1(_04351_),
    .X(_04438_));
 sky130_fd_sc_hd__xor2_1 _24262_ (.A(_04278_),
    .B(_04438_),
    .X(_04439_));
 sky130_fd_sc_hd__nand2_1 _24263_ (.A(_04363_),
    .B(_04439_),
    .Y(_04440_));
 sky130_fd_sc_hd__or2_1 _24264_ (.A(_04359_),
    .B(_04439_),
    .X(_04441_));
 sky130_fd_sc_hd__nand2_1 _24265_ (.A(_04440_),
    .B(_04441_),
    .Y(_04442_));
 sky130_fd_sc_hd__xor2_1 _24266_ (.A(_04437_),
    .B(_04442_),
    .X(_04443_));
 sky130_fd_sc_hd__or2_1 _24267_ (.A(_04355_),
    .B(_04357_),
    .X(_04444_));
 sky130_fd_sc_hd__o21a_1 _24268_ (.A1(_04358_),
    .A2(_04365_),
    .B1(_04444_),
    .X(_04445_));
 sky130_fd_sc_hd__xor2_1 _24269_ (.A(_04443_),
    .B(_04445_),
    .X(_04446_));
 sky130_fd_sc_hd__clkbuf_2 _24270_ (.A(_04278_),
    .X(_04447_));
 sky130_fd_sc_hd__a21oi_1 _24271_ (.A1(_04447_),
    .A2(_04360_),
    .B1(_04362_),
    .Y(_04448_));
 sky130_fd_sc_hd__xnor2_1 _24272_ (.A(_04208_),
    .B(_04448_),
    .Y(_04449_));
 sky130_fd_sc_hd__or2_1 _24273_ (.A(_04287_),
    .B(_04449_),
    .X(_04450_));
 sky130_fd_sc_hd__nand2_1 _24274_ (.A(_04287_),
    .B(_04449_),
    .Y(_04451_));
 sky130_fd_sc_hd__nand2_1 _24275_ (.A(_04450_),
    .B(_04451_),
    .Y(_04452_));
 sky130_fd_sc_hd__nor2_1 _24276_ (.A(_04446_),
    .B(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__and2_1 _24277_ (.A(_04446_),
    .B(_04452_),
    .X(_04454_));
 sky130_fd_sc_hd__nor2_1 _24278_ (.A(_04453_),
    .B(_04454_),
    .Y(_04455_));
 sky130_fd_sc_hd__o21ba_1 _24279_ (.A1(_04366_),
    .A2(_04368_),
    .B1_N(_04375_),
    .X(_04456_));
 sky130_fd_sc_hd__xnor2_1 _24280_ (.A(_04455_),
    .B(_04456_),
    .Y(_04457_));
 sky130_fd_sc_hd__clkbuf_2 _24281_ (.A(_04208_),
    .X(_04458_));
 sky130_fd_sc_hd__o21a_1 _24282_ (.A1(_04458_),
    .A2(_04370_),
    .B1(_04372_),
    .X(_04459_));
 sky130_fd_sc_hd__xnor2_1 _24283_ (.A(_04044_),
    .B(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hd__nor2_1 _24284_ (.A(_04222_),
    .B(_04460_),
    .Y(_04461_));
 sky130_fd_sc_hd__and2_1 _24285_ (.A(_04222_),
    .B(_04460_),
    .X(_04462_));
 sky130_fd_sc_hd__nor2_1 _24286_ (.A(_04461_),
    .B(_04462_),
    .Y(_04463_));
 sky130_fd_sc_hd__nand2_1 _24287_ (.A(_04457_),
    .B(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__or2_1 _24288_ (.A(_04457_),
    .B(_04463_),
    .X(_04465_));
 sky130_fd_sc_hd__nand2_1 _24289_ (.A(_04464_),
    .B(_04465_),
    .Y(_04466_));
 sky130_fd_sc_hd__o31a_1 _24290_ (.A1(_04375_),
    .A2(_04376_),
    .A3(_04378_),
    .B1(_04386_),
    .X(_04467_));
 sky130_fd_sc_hd__nor2_1 _24291_ (.A(_04466_),
    .B(_04467_),
    .Y(_04468_));
 sky130_fd_sc_hd__and2_1 _24292_ (.A(_04466_),
    .B(_04467_),
    .X(_04469_));
 sky130_fd_sc_hd__nor2_1 _24293_ (.A(_04468_),
    .B(_04469_),
    .Y(_04470_));
 sky130_fd_sc_hd__o21a_1 _24294_ (.A1(_04222_),
    .A2(_04384_),
    .B1(_04382_),
    .X(_04471_));
 sky130_fd_sc_hd__xnor2_1 _24295_ (.A(_03764_),
    .B(_04471_),
    .Y(_04472_));
 sky130_fd_sc_hd__nand2_1 _24296_ (.A(_04311_),
    .B(_04472_),
    .Y(_04473_));
 sky130_fd_sc_hd__or2_1 _24297_ (.A(_03874_),
    .B(_04472_),
    .X(_04474_));
 sky130_fd_sc_hd__and2_1 _24298_ (.A(_04473_),
    .B(_04474_),
    .X(_04475_));
 sky130_fd_sc_hd__xnor2_1 _24299_ (.A(_04470_),
    .B(_04475_),
    .Y(_04476_));
 sky130_fd_sc_hd__a21oi_1 _24300_ (.A1(_04392_),
    .A2(_04397_),
    .B1(_04390_),
    .Y(_04477_));
 sky130_fd_sc_hd__nor2_1 _24301_ (.A(_04476_),
    .B(_04477_),
    .Y(_04478_));
 sky130_fd_sc_hd__and2_1 _24302_ (.A(_04476_),
    .B(_04477_),
    .X(_04479_));
 sky130_fd_sc_hd__or2_1 _24303_ (.A(_04478_),
    .B(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__or3_1 _24304_ (.A(_04322_),
    .B(_04323_),
    .C(_04393_),
    .X(_04481_));
 sky130_fd_sc_hd__buf_1 _24305_ (.A(_04158_),
    .X(_04482_));
 sky130_fd_sc_hd__a21oi_1 _24306_ (.A1(_04481_),
    .A2(_04395_),
    .B1(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__and3_1 _24307_ (.A(_04482_),
    .B(_04481_),
    .C(_04395_),
    .X(_04484_));
 sky130_fd_sc_hd__or2_1 _24308_ (.A(_04483_),
    .B(_04484_),
    .X(_04485_));
 sky130_fd_sc_hd__nor2_1 _24309_ (.A(_04480_),
    .B(_04485_),
    .Y(_04486_));
 sky130_fd_sc_hd__and2_1 _24310_ (.A(_04480_),
    .B(_04485_),
    .X(_04487_));
 sky130_fd_sc_hd__nor2_1 _24311_ (.A(_04486_),
    .B(_04487_),
    .Y(_04488_));
 sky130_fd_sc_hd__o21ba_1 _24312_ (.A1(_04398_),
    .A2(_04400_),
    .B1_N(_04406_),
    .X(_04489_));
 sky130_fd_sc_hd__xnor2_1 _24313_ (.A(_04488_),
    .B(_04489_),
    .Y(_04490_));
 sky130_fd_sc_hd__nand2_1 _24314_ (.A(_04403_),
    .B(_04490_),
    .Y(_04491_));
 sky130_fd_sc_hd__or2_1 _24315_ (.A(_04403_),
    .B(_04490_),
    .X(_04492_));
 sky130_fd_sc_hd__nand2_1 _24316_ (.A(_04491_),
    .B(_04492_),
    .Y(_04493_));
 sky130_fd_sc_hd__a21oi_1 _24317_ (.A1(_04418_),
    .A2(_04419_),
    .B1(_04493_),
    .Y(_04494_));
 sky130_fd_sc_hd__and3_1 _24318_ (.A(_04418_),
    .B(_04419_),
    .C(_04493_),
    .X(_04495_));
 sky130_fd_sc_hd__nor2_1 _24319_ (.A(_04494_),
    .B(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__nand2_1 _24320_ (.A(_04170_),
    .B(_04251_),
    .Y(_04497_));
 sky130_fd_sc_hd__a211o_1 _24321_ (.A1(_03982_),
    .A2(_04172_),
    .B1(_04173_),
    .C1(_04497_),
    .X(_04498_));
 sky130_fd_sc_hd__o21a_1 _24322_ (.A1(_04335_),
    .A2(_04415_),
    .B1(_04413_),
    .X(_04499_));
 sky130_fd_sc_hd__nor2_1 _24323_ (.A(_04339_),
    .B(_04499_),
    .Y(_04500_));
 sky130_fd_sc_hd__nor2_1 _24324_ (.A(_04336_),
    .B(_04415_),
    .Y(_04501_));
 sky130_fd_sc_hd__a211oi_2 _24325_ (.A1(_04498_),
    .A2(_04500_),
    .B1(_04501_),
    .C1(_04414_),
    .Y(_04502_));
 sky130_fd_sc_hd__xor2_1 _24326_ (.A(_04496_),
    .B(_04502_),
    .X(_00106_));
 sky130_fd_sc_hd__or3_1 _24327_ (.A(_04486_),
    .B(_04487_),
    .C(_04489_),
    .X(_04503_));
 sky130_fd_sc_hd__and2b_1 _24328_ (.A_N(_04445_),
    .B(_04443_),
    .X(_04504_));
 sky130_fd_sc_hd__or2b_1 _24329_ (.A(_04436_),
    .B_N(_04434_),
    .X(_04505_));
 sky130_fd_sc_hd__o21a_1 _24330_ (.A1(_04437_),
    .A2(_04442_),
    .B1(_04505_),
    .X(_04506_));
 sky130_vsdinv _24331_ (.A(_13805_),
    .Y(_04507_));
 sky130_fd_sc_hd__o2bb2a_1 _24332_ (.A1_N(_13818_),
    .A2_N(_04257_),
    .B1(_04507_),
    .B2(_04264_),
    .X(_04508_));
 sky130_fd_sc_hd__and4b_1 _24333_ (.A_N(_04264_),
    .B(_14023_),
    .C(_04257_),
    .D(_13805_),
    .X(_04509_));
 sky130_fd_sc_hd__nor2_1 _24334_ (.A(_04508_),
    .B(_04509_),
    .Y(_04510_));
 sky130_fd_sc_hd__buf_2 _24335_ (.A(_04084_),
    .X(_04511_));
 sky130_fd_sc_hd__nand2_1 _24336_ (.A(_04511_),
    .B(_14213_),
    .Y(_04512_));
 sky130_fd_sc_hd__xnor2_1 _24337_ (.A(_04510_),
    .B(_04512_),
    .Y(_04513_));
 sky130_fd_sc_hd__o21ba_1 _24338_ (.A1(_04421_),
    .A2(_04424_),
    .B1_N(_04422_),
    .X(_04514_));
 sky130_fd_sc_hd__xnor2_1 _24339_ (.A(_04513_),
    .B(_04514_),
    .Y(_04515_));
 sky130_fd_sc_hd__or2_1 _24340_ (.A(_04094_),
    .B(_04091_),
    .X(_04516_));
 sky130_fd_sc_hd__and3b_1 _24341_ (.A_N(_04429_),
    .B(_04516_),
    .C(_14564_),
    .X(_04517_));
 sky130_fd_sc_hd__xnor2_2 _24342_ (.A(_04353_),
    .B(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__xnor2_1 _24343_ (.A(_04515_),
    .B(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__or2b_1 _24344_ (.A(_04425_),
    .B_N(_04426_),
    .X(_04520_));
 sky130_fd_sc_hd__and2b_1 _24345_ (.A_N(_04426_),
    .B(_04425_),
    .X(_04521_));
 sky130_fd_sc_hd__a21oi_1 _24346_ (.A1(_04520_),
    .A2(_04433_),
    .B1(_04521_),
    .Y(_04522_));
 sky130_fd_sc_hd__xnor2_1 _24347_ (.A(_04519_),
    .B(_04522_),
    .Y(_04523_));
 sky130_fd_sc_hd__o21a_1 _24348_ (.A1(_04430_),
    .A2(_04431_),
    .B1(_04447_),
    .X(_04524_));
 sky130_fd_sc_hd__nor3_1 _24349_ (.A(_04447_),
    .B(_04430_),
    .C(_04431_),
    .Y(_04525_));
 sky130_fd_sc_hd__nor2_1 _24350_ (.A(_04524_),
    .B(_04525_),
    .Y(_04526_));
 sky130_fd_sc_hd__xnor2_1 _24351_ (.A(_04363_),
    .B(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__xor2_1 _24352_ (.A(_04523_),
    .B(_04527_),
    .X(_04528_));
 sky130_fd_sc_hd__or2b_1 _24353_ (.A(_04506_),
    .B_N(_04528_),
    .X(_04529_));
 sky130_fd_sc_hd__or2b_1 _24354_ (.A(_04528_),
    .B_N(_04506_),
    .X(_04530_));
 sky130_fd_sc_hd__nand2_1 _24355_ (.A(_04529_),
    .B(_04530_),
    .Y(_04531_));
 sky130_fd_sc_hd__nand2_1 _24356_ (.A(_04447_),
    .B(_04438_),
    .Y(_04532_));
 sky130_fd_sc_hd__a21o_1 _24357_ (.A1(_04532_),
    .A2(_04440_),
    .B1(_04208_),
    .X(_04533_));
 sky130_fd_sc_hd__nand3_1 _24358_ (.A(_04458_),
    .B(_04532_),
    .C(_04440_),
    .Y(_04534_));
 sky130_fd_sc_hd__nand2_1 _24359_ (.A(_04533_),
    .B(_04534_),
    .Y(_04535_));
 sky130_fd_sc_hd__xnor2_1 _24360_ (.A(_04299_),
    .B(_04535_),
    .Y(_04536_));
 sky130_fd_sc_hd__xor2_1 _24361_ (.A(_04531_),
    .B(_04536_),
    .X(_04537_));
 sky130_fd_sc_hd__o21a_1 _24362_ (.A1(_04504_),
    .A2(_04453_),
    .B1(_04537_),
    .X(_04538_));
 sky130_fd_sc_hd__nor3_1 _24363_ (.A(_04504_),
    .B(_04453_),
    .C(_04537_),
    .Y(_04539_));
 sky130_fd_sc_hd__nor2_1 _24364_ (.A(_04538_),
    .B(_04539_),
    .Y(_04540_));
 sky130_fd_sc_hd__o21a_1 _24365_ (.A1(_04458_),
    .A2(_04448_),
    .B1(_04450_),
    .X(_04541_));
 sky130_fd_sc_hd__xnor2_1 _24366_ (.A(_04229_),
    .B(_04541_),
    .Y(_04542_));
 sky130_fd_sc_hd__nor2_1 _24367_ (.A(_04298_),
    .B(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hd__and2_1 _24368_ (.A(_04222_),
    .B(_04542_),
    .X(_04544_));
 sky130_fd_sc_hd__nor2_1 _24369_ (.A(_04543_),
    .B(_04544_),
    .Y(_04545_));
 sky130_fd_sc_hd__xnor2_1 _24370_ (.A(_04540_),
    .B(_04545_),
    .Y(_04546_));
 sky130_fd_sc_hd__o31a_1 _24371_ (.A1(_04453_),
    .A2(_04454_),
    .A3(_04456_),
    .B1(_04464_),
    .X(_04547_));
 sky130_fd_sc_hd__nor2_1 _24372_ (.A(_04546_),
    .B(_04547_),
    .Y(_04548_));
 sky130_fd_sc_hd__and2_1 _24373_ (.A(_04546_),
    .B(_04547_),
    .X(_04549_));
 sky130_fd_sc_hd__nor2_1 _24374_ (.A(_04548_),
    .B(_04549_),
    .Y(_04550_));
 sky130_fd_sc_hd__o21ba_1 _24375_ (.A1(_04312_),
    .A2(_04459_),
    .B1_N(_04461_),
    .X(_04551_));
 sky130_fd_sc_hd__xnor2_1 _24376_ (.A(_04156_),
    .B(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__nand2_1 _24377_ (.A(_04311_),
    .B(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__or2_1 _24378_ (.A(_03874_),
    .B(_04552_),
    .X(_04554_));
 sky130_fd_sc_hd__and2_1 _24379_ (.A(_04553_),
    .B(_04554_),
    .X(_04555_));
 sky130_fd_sc_hd__xnor2_1 _24380_ (.A(_04550_),
    .B(_04555_),
    .Y(_04556_));
 sky130_fd_sc_hd__a21oi_1 _24381_ (.A1(_04470_),
    .A2(_04475_),
    .B1(_04468_),
    .Y(_04557_));
 sky130_fd_sc_hd__or2_1 _24382_ (.A(_04556_),
    .B(_04557_),
    .X(_04558_));
 sky130_fd_sc_hd__nand2_1 _24383_ (.A(_04556_),
    .B(_04557_),
    .Y(_04559_));
 sky130_fd_sc_hd__nand2_1 _24384_ (.A(_04558_),
    .B(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__or3_1 _24385_ (.A(_04322_),
    .B(_04323_),
    .C(_04471_),
    .X(_04561_));
 sky130_fd_sc_hd__a21oi_1 _24386_ (.A1(_04561_),
    .A2(_04473_),
    .B1(_04482_),
    .Y(_04562_));
 sky130_fd_sc_hd__and3_1 _24387_ (.A(_04482_),
    .B(_04561_),
    .C(_04473_),
    .X(_04563_));
 sky130_fd_sc_hd__or2_1 _24388_ (.A(_04562_),
    .B(_04563_),
    .X(_04564_));
 sky130_fd_sc_hd__xor2_1 _24389_ (.A(_04560_),
    .B(_04564_),
    .X(_04565_));
 sky130_fd_sc_hd__o21ai_1 _24390_ (.A1(_04478_),
    .A2(_04486_),
    .B1(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hd__or3_1 _24391_ (.A(_04478_),
    .B(_04486_),
    .C(_04565_),
    .X(_04567_));
 sky130_fd_sc_hd__and2_1 _24392_ (.A(_04566_),
    .B(_04567_),
    .X(_04568_));
 sky130_fd_sc_hd__nand2_1 _24393_ (.A(_04483_),
    .B(_04568_),
    .Y(_04569_));
 sky130_fd_sc_hd__or2_1 _24394_ (.A(_04483_),
    .B(_04568_),
    .X(_04570_));
 sky130_fd_sc_hd__nand2_1 _24395_ (.A(_04569_),
    .B(_04570_),
    .Y(_04571_));
 sky130_fd_sc_hd__a21oi_1 _24396_ (.A1(_04503_),
    .A2(_04491_),
    .B1(_04571_),
    .Y(_04572_));
 sky130_fd_sc_hd__nand3_1 _24397_ (.A(_04503_),
    .B(_04491_),
    .C(_04571_),
    .Y(_04573_));
 sky130_fd_sc_hd__or2b_1 _24398_ (.A(_04572_),
    .B_N(_04573_),
    .X(_04574_));
 sky130_fd_sc_hd__a21o_1 _24399_ (.A1(_04496_),
    .A2(_04502_),
    .B1(_04494_),
    .X(_04575_));
 sky130_fd_sc_hd__xnor2_1 _24400_ (.A(_04574_),
    .B(_04575_),
    .Y(_00107_));
 sky130_fd_sc_hd__o21a_1 _24401_ (.A1(_04560_),
    .A2(_04564_),
    .B1(_04558_),
    .X(_04576_));
 sky130_fd_sc_hd__o21a_1 _24402_ (.A1(_04531_),
    .A2(_04536_),
    .B1(_04529_),
    .X(_04577_));
 sky130_fd_sc_hd__or2_1 _24403_ (.A(_04519_),
    .B(_04522_),
    .X(_04578_));
 sky130_fd_sc_hd__o21a_1 _24404_ (.A1(_04523_),
    .A2(_04527_),
    .B1(_04578_),
    .X(_04579_));
 sky130_fd_sc_hd__or2b_1 _24405_ (.A(_04514_),
    .B_N(_04513_),
    .X(_04580_));
 sky130_fd_sc_hd__nand2_1 _24406_ (.A(_04515_),
    .B(_04518_),
    .Y(_04581_));
 sky130_fd_sc_hd__and3_1 _24407_ (.A(_04511_),
    .B(_14214_),
    .C(_04510_),
    .X(_04582_));
 sky130_fd_sc_hd__nor2_1 _24408_ (.A(_13819_),
    .B(_04507_),
    .Y(_04583_));
 sky130_fd_sc_hd__and2_1 _24409_ (.A(_04254_),
    .B(_03628_),
    .X(_04584_));
 sky130_fd_sc_hd__nor2_1 _24410_ (.A(_04583_),
    .B(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__and2_1 _24411_ (.A(_04583_),
    .B(_04584_),
    .X(_04586_));
 sky130_fd_sc_hd__nor2_1 _24412_ (.A(_04585_),
    .B(_04586_),
    .Y(_04587_));
 sky130_fd_sc_hd__nand2_1 _24413_ (.A(_04511_),
    .B(_14565_),
    .Y(_04588_));
 sky130_fd_sc_hd__xnor2_1 _24414_ (.A(_04587_),
    .B(_04588_),
    .Y(_04589_));
 sky130_fd_sc_hd__o21ai_1 _24415_ (.A1(_04509_),
    .A2(_04582_),
    .B1(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__or3_1 _24416_ (.A(_04509_),
    .B(_04582_),
    .C(_04589_),
    .X(_04591_));
 sky130_fd_sc_hd__nand2_1 _24417_ (.A(_04590_),
    .B(_04591_),
    .Y(_04592_));
 sky130_fd_sc_hd__xor2_1 _24418_ (.A(_04518_),
    .B(_04592_),
    .X(_04593_));
 sky130_fd_sc_hd__a21o_1 _24419_ (.A1(_04580_),
    .A2(_04581_),
    .B1(_04593_),
    .X(_04594_));
 sky130_fd_sc_hd__nand3_1 _24420_ (.A(_04580_),
    .B(_04581_),
    .C(_04593_),
    .Y(_04595_));
 sky130_fd_sc_hd__nand2_1 _24421_ (.A(_04594_),
    .B(_04595_),
    .Y(_04596_));
 sky130_fd_sc_hd__a31o_1 _24422_ (.A1(_04098_),
    .A2(_14565_),
    .A3(_04516_),
    .B1(_04429_),
    .X(_04597_));
 sky130_fd_sc_hd__xor2_1 _24423_ (.A(_04447_),
    .B(_04597_),
    .X(_04598_));
 sky130_fd_sc_hd__and2_1 _24424_ (.A(_04363_),
    .B(_04598_),
    .X(_04599_));
 sky130_fd_sc_hd__nor2_1 _24425_ (.A(_04363_),
    .B(_04598_),
    .Y(_04600_));
 sky130_fd_sc_hd__or2_1 _24426_ (.A(_04599_),
    .B(_04600_),
    .X(_04601_));
 sky130_fd_sc_hd__xnor2_1 _24427_ (.A(_04596_),
    .B(_04601_),
    .Y(_04602_));
 sky130_fd_sc_hd__xnor2_1 _24428_ (.A(_04579_),
    .B(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__a21oi_1 _24429_ (.A1(_04363_),
    .A2(_04526_),
    .B1(_04524_),
    .Y(_04604_));
 sky130_fd_sc_hd__xnor2_1 _24430_ (.A(_04458_),
    .B(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__xnor2_1 _24431_ (.A(_04299_),
    .B(_04605_),
    .Y(_04606_));
 sky130_fd_sc_hd__or2_1 _24432_ (.A(_04603_),
    .B(_04606_),
    .X(_04607_));
 sky130_fd_sc_hd__nand2_1 _24433_ (.A(_04603_),
    .B(_04606_),
    .Y(_04608_));
 sky130_fd_sc_hd__and2_1 _24434_ (.A(_04607_),
    .B(_04608_),
    .X(_04609_));
 sky130_fd_sc_hd__and2b_1 _24435_ (.A_N(_04577_),
    .B(_04609_),
    .X(_04610_));
 sky130_fd_sc_hd__and2b_1 _24436_ (.A_N(_04609_),
    .B(_04577_),
    .X(_04611_));
 sky130_fd_sc_hd__or2_1 _24437_ (.A(_04610_),
    .B(_04611_),
    .X(_04612_));
 sky130_fd_sc_hd__o21a_1 _24438_ (.A1(_04299_),
    .A2(_04535_),
    .B1(_04533_),
    .X(_04613_));
 sky130_fd_sc_hd__or2_1 _24439_ (.A(_04312_),
    .B(_04613_),
    .X(_04614_));
 sky130_fd_sc_hd__nand2_1 _24440_ (.A(_04312_),
    .B(_04613_),
    .Y(_04615_));
 sky130_fd_sc_hd__nand2_1 _24441_ (.A(_04614_),
    .B(_04615_),
    .Y(_04616_));
 sky130_fd_sc_hd__xor2_1 _24442_ (.A(_04298_),
    .B(_04616_),
    .X(_04617_));
 sky130_fd_sc_hd__xor2_1 _24443_ (.A(_04612_),
    .B(_04617_),
    .X(_04618_));
 sky130_fd_sc_hd__a21oi_1 _24444_ (.A1(_04540_),
    .A2(_04545_),
    .B1(_04538_),
    .Y(_04619_));
 sky130_fd_sc_hd__xnor2_1 _24445_ (.A(_04618_),
    .B(_04619_),
    .Y(_04620_));
 sky130_fd_sc_hd__o21ba_1 _24446_ (.A1(_04312_),
    .A2(_04541_),
    .B1_N(_04543_),
    .X(_04621_));
 sky130_fd_sc_hd__xnor2_1 _24447_ (.A(_04156_),
    .B(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__nand2_1 _24448_ (.A(_04311_),
    .B(_04622_),
    .Y(_04623_));
 sky130_fd_sc_hd__or2_1 _24449_ (.A(_04311_),
    .B(_04622_),
    .X(_04624_));
 sky130_fd_sc_hd__and2_1 _24450_ (.A(_04623_),
    .B(_04624_),
    .X(_04625_));
 sky130_fd_sc_hd__xor2_1 _24451_ (.A(_04620_),
    .B(_04625_),
    .X(_04626_));
 sky130_fd_sc_hd__a21oi_1 _24452_ (.A1(_04550_),
    .A2(_04555_),
    .B1(_04548_),
    .Y(_04627_));
 sky130_fd_sc_hd__or2_1 _24453_ (.A(_04626_),
    .B(_04627_),
    .X(_04628_));
 sky130_fd_sc_hd__nand2_1 _24454_ (.A(_04626_),
    .B(_04627_),
    .Y(_04629_));
 sky130_fd_sc_hd__nand2_1 _24455_ (.A(_04628_),
    .B(_04629_),
    .Y(_04630_));
 sky130_fd_sc_hd__o31a_1 _24456_ (.A1(_04322_),
    .A2(_04323_),
    .A3(_04551_),
    .B1(_04553_),
    .X(_04631_));
 sky130_fd_sc_hd__and2b_1 _24457_ (.A_N(_04482_),
    .B(_04631_),
    .X(_04632_));
 sky130_fd_sc_hd__and2b_1 _24458_ (.A_N(_04631_),
    .B(_04482_),
    .X(_04633_));
 sky130_fd_sc_hd__nor2_1 _24459_ (.A(_04632_),
    .B(_04633_),
    .Y(_04634_));
 sky130_fd_sc_hd__xor2_1 _24460_ (.A(_04630_),
    .B(_04634_),
    .X(_04635_));
 sky130_fd_sc_hd__and2b_1 _24461_ (.A_N(_04576_),
    .B(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__and2b_1 _24462_ (.A_N(_04635_),
    .B(_04576_),
    .X(_04637_));
 sky130_fd_sc_hd__nor2_1 _24463_ (.A(_04636_),
    .B(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__xnor2_1 _24464_ (.A(_04562_),
    .B(_04638_),
    .Y(_04639_));
 sky130_fd_sc_hd__a21o_1 _24465_ (.A1(_04566_),
    .A2(_04569_),
    .B1(_04639_),
    .X(_04640_));
 sky130_fd_sc_hd__nand3_1 _24466_ (.A(_04566_),
    .B(_04569_),
    .C(_04639_),
    .Y(_04641_));
 sky130_fd_sc_hd__nand2_1 _24467_ (.A(_04640_),
    .B(_04641_),
    .Y(_04642_));
 sky130_fd_sc_hd__and2_1 _24468_ (.A(_04494_),
    .B(_04573_),
    .X(_04643_));
 sky130_fd_sc_hd__a311o_1 _24469_ (.A1(_04496_),
    .A2(_04502_),
    .A3(_04573_),
    .B1(_04643_),
    .C1(_04572_),
    .X(_04644_));
 sky130_fd_sc_hd__xnor2_1 _24470_ (.A(_04642_),
    .B(_04644_),
    .Y(_00108_));
 sky130_fd_sc_hd__a21bo_1 _24471_ (.A1(_04641_),
    .A2(_04644_),
    .B1_N(_04640_),
    .X(_04645_));
 sky130_fd_sc_hd__a21oi_1 _24472_ (.A1(_04562_),
    .A2(_04638_),
    .B1(_04636_),
    .Y(_04646_));
 sky130_fd_sc_hd__o21ai_1 _24473_ (.A1(_04630_),
    .A2(_04634_),
    .B1(_04628_),
    .Y(_04647_));
 sky130_fd_sc_hd__or2b_1 _24474_ (.A(_04620_),
    .B_N(_04625_),
    .X(_04648_));
 sky130_fd_sc_hd__o21a_1 _24475_ (.A1(_04618_),
    .A2(_04619_),
    .B1(_04648_),
    .X(_04649_));
 sky130_vsdinv _24476_ (.A(_04612_),
    .Y(_04650_));
 sky130_fd_sc_hd__a21o_1 _24477_ (.A1(_04650_),
    .A2(_04617_),
    .B1(_04610_),
    .X(_04651_));
 sky130_fd_sc_hd__o21ai_1 _24478_ (.A1(_04579_),
    .A2(_04602_),
    .B1(_04607_),
    .Y(_04652_));
 sky130_fd_sc_hd__or2_1 _24479_ (.A(_04458_),
    .B(_04604_),
    .X(_04653_));
 sky130_fd_sc_hd__o21ai_1 _24480_ (.A1(_04299_),
    .A2(_04605_),
    .B1(_04653_),
    .Y(_04654_));
 sky130_fd_sc_hd__mux2_1 _24481_ (.A0(_04595_),
    .A1(_04594_),
    .S(_04601_),
    .X(_04655_));
 sky130_fd_sc_hd__xnor2_1 _24482_ (.A(_04654_),
    .B(_04655_),
    .Y(_04656_));
 sky130_fd_sc_hd__mux2_1 _24483_ (.A0(_04590_),
    .A1(_04591_),
    .S(_04518_),
    .X(_04657_));
 sky130_fd_sc_hd__o21ba_1 _24484_ (.A1(_04585_),
    .A2(_04588_),
    .B1_N(_04586_),
    .X(_04658_));
 sky130_fd_sc_hd__nor2_1 _24485_ (.A(_14214_),
    .B(_04507_),
    .Y(_04659_));
 sky130_fd_sc_hd__o21ai_1 _24486_ (.A1(_04511_),
    .A2(_04254_),
    .B1(_14565_),
    .Y(_04660_));
 sky130_fd_sc_hd__a21oi_1 _24487_ (.A1(_04511_),
    .A2(_04254_),
    .B1(_04660_),
    .Y(_04661_));
 sky130_fd_sc_hd__xnor2_1 _24488_ (.A(_04659_),
    .B(_04661_),
    .Y(_04662_));
 sky130_fd_sc_hd__xnor2_1 _24489_ (.A(_04658_),
    .B(_04662_),
    .Y(_04663_));
 sky130_fd_sc_hd__xnor2_1 _24490_ (.A(_04657_),
    .B(_04663_),
    .Y(_04664_));
 sky130_fd_sc_hd__a21oi_1 _24491_ (.A1(_04447_),
    .A2(_04597_),
    .B1(_04599_),
    .Y(_04665_));
 sky130_fd_sc_hd__mux2_1 _24492_ (.A0(_04120_),
    .A1(_04299_),
    .S(_04458_),
    .X(_04666_));
 sky130_fd_sc_hd__xnor2_1 _24493_ (.A(_04665_),
    .B(_04666_),
    .Y(_04667_));
 sky130_fd_sc_hd__xnor2_1 _24494_ (.A(_04664_),
    .B(_04667_),
    .Y(_04668_));
 sky130_fd_sc_hd__mux2_1 _24495_ (.A0(_03948_),
    .A1(_04298_),
    .S(_04312_),
    .X(_04669_));
 sky130_fd_sc_hd__xnor2_1 _24496_ (.A(_04668_),
    .B(_04669_),
    .Y(_04670_));
 sky130_fd_sc_hd__xnor2_1 _24497_ (.A(_04656_),
    .B(_04670_),
    .Y(_04671_));
 sky130_fd_sc_hd__xnor2_1 _24498_ (.A(_04652_),
    .B(_04671_),
    .Y(_04672_));
 sky130_fd_sc_hd__mux2_1 _24499_ (.A0(_03478_),
    .A1(_03361_),
    .S(_04156_),
    .X(_04673_));
 sky130_fd_sc_hd__o21ai_1 _24500_ (.A1(_04298_),
    .A2(_04616_),
    .B1(_04614_),
    .Y(_04674_));
 sky130_fd_sc_hd__xnor2_1 _24501_ (.A(_04673_),
    .B(_04674_),
    .Y(_04675_));
 sky130_fd_sc_hd__xnor2_1 _24502_ (.A(_04672_),
    .B(_04675_),
    .Y(_04676_));
 sky130_fd_sc_hd__xnor2_1 _24503_ (.A(_04651_),
    .B(_04676_),
    .Y(_04677_));
 sky130_fd_sc_hd__o31a_1 _24504_ (.A1(_04322_),
    .A2(_04323_),
    .A3(_04621_),
    .B1(_04623_),
    .X(_04678_));
 sky130_fd_sc_hd__xnor2_1 _24505_ (.A(_04632_),
    .B(_04678_),
    .Y(_04679_));
 sky130_fd_sc_hd__xnor2_1 _24506_ (.A(_04677_),
    .B(_04679_),
    .Y(_04680_));
 sky130_fd_sc_hd__xnor2_1 _24507_ (.A(_04649_),
    .B(_04680_),
    .Y(_04681_));
 sky130_fd_sc_hd__xnor2_1 _24508_ (.A(_04647_),
    .B(_04681_),
    .Y(_04682_));
 sky130_fd_sc_hd__xnor2_1 _24509_ (.A(_04646_),
    .B(_04682_),
    .Y(_04683_));
 sky130_fd_sc_hd__xnor2_1 _24510_ (.A(_04645_),
    .B(_04683_),
    .Y(_00109_));
 sky130_fd_sc_hd__nor2_1 _24511_ (.A(_10690_),
    .B(_10733_),
    .Y(_04684_));
 sky130_fd_sc_hd__o32a_1 _24512_ (.A1(_10620_),
    .A2(_10658_),
    .A3(_10692_),
    .B1(_10777_),
    .B2(_04684_),
    .X(_04685_));
 sky130_fd_sc_hd__nor2_1 _24513_ (.A(_10734_),
    .B(_04685_),
    .Y(_00055_));
 sky130_fd_sc_hd__buf_2 _24514_ (.A(net161),
    .X(_04686_));
 sky130_fd_sc_hd__mux2_1 _24515_ (.A0(_08482_),
    .A1(_08460_),
    .S(_04686_),
    .X(_04687_));
 sky130_fd_sc_hd__mux2_1 _24516_ (.A0(_08407_),
    .A1(_08449_),
    .S(_08469_),
    .X(_04688_));
 sky130_fd_sc_hd__mux2_1 _24517_ (.A0(_04687_),
    .A1(_04688_),
    .S(_10105_),
    .X(_04689_));
 sky130_fd_sc_hd__mux2_1 _24518_ (.A0(_08475_),
    .A1(_08441_),
    .S(_04686_),
    .X(_04690_));
 sky130_fd_sc_hd__mux2_1 _24519_ (.A0(_08456_),
    .A1(_08679_),
    .S(_04686_),
    .X(_04691_));
 sky130_fd_sc_hd__buf_2 _24520_ (.A(net172),
    .X(_04692_));
 sky130_fd_sc_hd__mux2_1 _24521_ (.A0(_04690_),
    .A1(_04691_),
    .S(_04692_),
    .X(_04693_));
 sky130_fd_sc_hd__buf_2 _24522_ (.A(_08455_),
    .X(_04694_));
 sky130_fd_sc_hd__mux2_1 _24523_ (.A0(_04689_),
    .A1(_04693_),
    .S(_04694_),
    .X(_04695_));
 sky130_fd_sc_hd__buf_2 _24524_ (.A(net161),
    .X(_04696_));
 sky130_fd_sc_hd__mux2_1 _24525_ (.A0(_08378_),
    .A1(_10186_),
    .S(_04696_),
    .X(_04697_));
 sky130_fd_sc_hd__mux2_1 _24526_ (.A0(_08417_),
    .A1(_08346_),
    .S(_04696_),
    .X(_04698_));
 sky130_fd_sc_hd__mux2_1 _24527_ (.A0(_08342_),
    .A1(_08411_),
    .S(_04686_),
    .X(_04699_));
 sky130_fd_sc_hd__mux2_1 _24528_ (.A0(_08401_),
    .A1(_10156_),
    .S(_04686_),
    .X(_04700_));
 sky130_fd_sc_hd__clkbuf_2 _24529_ (.A(_10271_),
    .X(_04701_));
 sky130_fd_sc_hd__mux4_1 _24530_ (.A0(_04697_),
    .A1(_04698_),
    .A2(_04699_),
    .A3(_04700_),
    .S0(_10284_),
    .S1(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__mux2_1 _24531_ (.A0(_04695_),
    .A1(_04702_),
    .S(_10431_),
    .X(_04703_));
 sky130_fd_sc_hd__buf_2 _24532_ (.A(_08443_),
    .X(_04704_));
 sky130_fd_sc_hd__clkbuf_2 _24533_ (.A(_04704_),
    .X(_04705_));
 sky130_fd_sc_hd__clkbuf_2 _24534_ (.A(_08455_),
    .X(_04706_));
 sky130_fd_sc_hd__nand2_1 _24535_ (.A(_08325_),
    .B(_08470_),
    .Y(_04707_));
 sky130_fd_sc_hd__or3_1 _24536_ (.A(_10285_),
    .B(_04706_),
    .C(_04707_),
    .X(_04708_));
 sky130_fd_sc_hd__nor2_1 _24537_ (.A(_04705_),
    .B(_04708_),
    .Y(_04709_));
 sky130_fd_sc_hd__buf_2 _24538_ (.A(_10276_),
    .X(_04710_));
 sky130_fd_sc_hd__mux2_1 _24539_ (.A0(_04703_),
    .A1(_04709_),
    .S(_04710_),
    .X(_04711_));
 sky130_fd_sc_hd__clkbuf_1 _24540_ (.A(_04711_),
    .X(_14604_));
 sky130_fd_sc_hd__buf_2 _24541_ (.A(_10105_),
    .X(_04712_));
 sky130_fd_sc_hd__mux4_1 _24542_ (.A0(_10156_),
    .A1(_08482_),
    .A2(_08460_),
    .A3(_10337_),
    .S0(_10268_),
    .S1(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__mux4_1 _24543_ (.A0(_10334_),
    .A1(_08475_),
    .A2(_08441_),
    .A3(_08456_),
    .S0(_10268_),
    .S1(_04712_),
    .X(_04714_));
 sky130_fd_sc_hd__mux2_1 _24544_ (.A0(_04713_),
    .A1(_04714_),
    .S(_04694_),
    .X(_04715_));
 sky130_fd_sc_hd__clkbuf_2 _24545_ (.A(_10105_),
    .X(_04716_));
 sky130_fd_sc_hd__mux4_1 _24546_ (.A0(_10197_),
    .A1(_08378_),
    .A2(_10186_),
    .A3(_10361_),
    .S0(_10281_),
    .S1(_04716_),
    .X(_04717_));
 sky130_fd_sc_hd__buf_2 _24547_ (.A(_08469_),
    .X(_04718_));
 sky130_fd_sc_hd__mux4_1 _24548_ (.A0(_08346_),
    .A1(_08342_),
    .A2(_08411_),
    .A3(_08401_),
    .S0(_04718_),
    .S1(_04712_),
    .X(_04719_));
 sky130_fd_sc_hd__mux2_1 _24549_ (.A0(_04717_),
    .A1(_04719_),
    .S(_04694_),
    .X(_04720_));
 sky130_fd_sc_hd__mux2_1 _24550_ (.A0(_04715_),
    .A1(_04720_),
    .S(_10431_),
    .X(_04721_));
 sky130_fd_sc_hd__clkbuf_2 _24551_ (.A(_08455_),
    .X(_04722_));
 sky130_fd_sc_hd__clkbuf_2 _24552_ (.A(_04722_),
    .X(_04723_));
 sky130_fd_sc_hd__a21oi_1 _24553_ (.A1(_08758_),
    .A2(_08470_),
    .B1(_08471_),
    .Y(_04724_));
 sky130_fd_sc_hd__or2_1 _24554_ (.A(_10106_),
    .B(_04724_),
    .X(_04725_));
 sky130_fd_sc_hd__or2_1 _24555_ (.A(_04723_),
    .B(_04725_),
    .X(_04726_));
 sky130_fd_sc_hd__nor2_1 _24556_ (.A(_04705_),
    .B(_04726_),
    .Y(_04727_));
 sky130_fd_sc_hd__mux2_1 _24557_ (.A0(_04721_),
    .A1(_04727_),
    .S(_04710_),
    .X(_04728_));
 sky130_fd_sc_hd__clkbuf_1 _24558_ (.A(_04728_),
    .X(_14605_));
 sky130_fd_sc_hd__mux2_1 _24559_ (.A0(_08351_),
    .A1(_08382_),
    .S(_04696_),
    .X(_04729_));
 sky130_fd_sc_hd__mux2_1 _24560_ (.A0(_04729_),
    .A1(_04697_),
    .S(_04712_),
    .X(_04730_));
 sky130_fd_sc_hd__mux2_1 _24561_ (.A0(_04698_),
    .A1(_04699_),
    .S(_04692_),
    .X(_04731_));
 sky130_fd_sc_hd__mux2_1 _24562_ (.A0(_04730_),
    .A1(_04731_),
    .S(_04701_),
    .X(_04732_));
 sky130_fd_sc_hd__mux2_1 _24563_ (.A0(_04700_),
    .A1(_04687_),
    .S(_04692_),
    .X(_04733_));
 sky130_fd_sc_hd__mux2_1 _24564_ (.A0(_04688_),
    .A1(_04690_),
    .S(_04692_),
    .X(_04734_));
 sky130_fd_sc_hd__mux2_1 _24565_ (.A0(_04733_),
    .A1(_04734_),
    .S(_04722_),
    .X(_04735_));
 sky130_fd_sc_hd__mux2_1 _24566_ (.A0(_04732_),
    .A1(_04735_),
    .S(_04704_),
    .X(_04736_));
 sky130_vsdinv _24567_ (.A(_04691_),
    .Y(_04737_));
 sky130_fd_sc_hd__mux2_1 _24568_ (.A0(_04737_),
    .A1(_04707_),
    .S(_10106_),
    .X(_04738_));
 sky130_fd_sc_hd__or2_1 _24569_ (.A(_10287_),
    .B(_04738_),
    .X(_04739_));
 sky130_fd_sc_hd__nor2_1 _24570_ (.A(_04705_),
    .B(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__mux2_1 _24571_ (.A0(_04736_),
    .A1(_04740_),
    .S(_04710_),
    .X(_04741_));
 sky130_fd_sc_hd__clkbuf_1 _24572_ (.A(_04741_),
    .X(_14606_));
 sky130_fd_sc_hd__mux4_1 _24573_ (.A0(_08411_),
    .A1(_08401_),
    .A2(_10156_),
    .A3(_10344_),
    .S0(_04718_),
    .S1(_04716_),
    .X(_04742_));
 sky130_fd_sc_hd__mux4_1 _24574_ (.A0(_08460_),
    .A1(_08407_),
    .A2(_08449_),
    .A3(_10331_),
    .S0(_10268_),
    .S1(_04712_),
    .X(_04743_));
 sky130_fd_sc_hd__mux2_1 _24575_ (.A0(_04742_),
    .A1(_04743_),
    .S(_04722_),
    .X(_04744_));
 sky130_fd_sc_hd__mux4_1 _24576_ (.A0(_10206_),
    .A1(_10372_),
    .A2(_08382_),
    .A3(_10367_),
    .S0(_10281_),
    .S1(_04716_),
    .X(_04745_));
 sky130_fd_sc_hd__mux4_1 _24577_ (.A0(_10186_),
    .A1(_08417_),
    .A2(_10357_),
    .A3(_08342_),
    .S0(_04718_),
    .S1(_04716_),
    .X(_04746_));
 sky130_fd_sc_hd__mux2_1 _24578_ (.A0(_04745_),
    .A1(_04746_),
    .S(_04694_),
    .X(_04747_));
 sky130_fd_sc_hd__mux2_1 _24579_ (.A0(_04744_),
    .A1(_04747_),
    .S(_10431_),
    .X(_04748_));
 sky130_fd_sc_hd__clkbuf_4 _24580_ (.A(_08469_),
    .X(_04749_));
 sky130_fd_sc_hd__mux4_2 _24581_ (.A0(_10322_),
    .A1(_10311_),
    .A2(_08758_),
    .A3(_08325_),
    .S0(_04749_),
    .S1(_10106_),
    .X(_04750_));
 sky130_fd_sc_hd__or2b_1 _24582_ (.A(_04723_),
    .B_N(_04750_),
    .X(_04751_));
 sky130_fd_sc_hd__nor2_1 _24583_ (.A(_04705_),
    .B(_04751_),
    .Y(_04752_));
 sky130_fd_sc_hd__buf_2 _24584_ (.A(_10276_),
    .X(_04753_));
 sky130_fd_sc_hd__mux2_1 _24585_ (.A0(_04748_),
    .A1(_04752_),
    .S(_04753_),
    .X(_04754_));
 sky130_fd_sc_hd__clkbuf_1 _24586_ (.A(_04754_),
    .X(_14607_));
 sky130_fd_sc_hd__clkbuf_4 _24587_ (.A(_10276_),
    .X(_04755_));
 sky130_fd_sc_hd__clkbuf_4 _24588_ (.A(_04755_),
    .X(_04756_));
 sky130_fd_sc_hd__buf_2 _24589_ (.A(_10271_),
    .X(_04757_));
 sky130_fd_sc_hd__buf_2 _24590_ (.A(_10284_),
    .X(_04758_));
 sky130_fd_sc_hd__o21ai_1 _24591_ (.A1(_04758_),
    .A2(_04707_),
    .B1(_10287_),
    .Y(_04759_));
 sky130_fd_sc_hd__o21ai_1 _24592_ (.A1(_04757_),
    .A2(_04693_),
    .B1(_04759_),
    .Y(_04760_));
 sky130_vsdinv _24593_ (.A(_04760_),
    .Y(_04761_));
 sky130_fd_sc_hd__clkbuf_2 _24594_ (.A(_10298_),
    .X(_04762_));
 sky130_fd_sc_hd__clkbuf_2 _24595_ (.A(_04762_),
    .X(_04763_));
 sky130_fd_sc_hd__buf_2 _24596_ (.A(_04692_),
    .X(_04764_));
 sky130_fd_sc_hd__mux2_1 _24597_ (.A0(_04699_),
    .A1(_04700_),
    .S(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__or2b_1 _24598_ (.A(_04689_),
    .B_N(_10272_),
    .X(_04766_));
 sky130_fd_sc_hd__o21ai_2 _24599_ (.A1(_04723_),
    .A2(_04765_),
    .B1(_04766_),
    .Y(_04767_));
 sky130_fd_sc_hd__buf_2 _24600_ (.A(_10298_),
    .X(_04768_));
 sky130_fd_sc_hd__mux2_1 _24601_ (.A0(_10378_),
    .A1(_08374_),
    .S(_04749_),
    .X(_04769_));
 sky130_fd_sc_hd__clkbuf_2 _24602_ (.A(_04722_),
    .X(_04770_));
 sky130_fd_sc_hd__mux4_1 _24603_ (.A0(_04769_),
    .A1(_04729_),
    .A2(_04697_),
    .A3(_04698_),
    .S0(_10107_),
    .S1(_04770_),
    .X(_04771_));
 sky130_fd_sc_hd__nor2_1 _24604_ (.A(_04768_),
    .B(_04771_),
    .Y(_04772_));
 sky130_fd_sc_hd__clkbuf_2 _24605_ (.A(_10276_),
    .X(_04773_));
 sky130_fd_sc_hd__a211oi_1 _24606_ (.A1(_04763_),
    .A2(_04767_),
    .B1(_04772_),
    .C1(_04773_),
    .Y(_04774_));
 sky130_fd_sc_hd__a31o_1 _24607_ (.A1(_10431_),
    .A2(_04756_),
    .A3(_04761_),
    .B1(_04774_),
    .X(_14608_));
 sky130_fd_sc_hd__mux4_1 _24608_ (.A0(_10214_),
    .A1(_10378_),
    .A2(_08374_),
    .A3(_10372_),
    .S0(_04749_),
    .S1(_04716_),
    .X(_04775_));
 sky130_fd_sc_hd__mux2_1 _24609_ (.A0(_04775_),
    .A1(_04717_),
    .S(_04701_),
    .X(_04776_));
 sky130_fd_sc_hd__mux2_1 _24610_ (.A0(_04719_),
    .A1(_04713_),
    .S(_04722_),
    .X(_04777_));
 sky130_fd_sc_hd__mux2_1 _24611_ (.A0(_04776_),
    .A1(_04777_),
    .S(_04704_),
    .X(_04778_));
 sky130_vsdinv _24612_ (.A(_04714_),
    .Y(_04779_));
 sky130_fd_sc_hd__mux2_1 _24613_ (.A0(_04779_),
    .A1(_04725_),
    .S(_04706_),
    .X(_04780_));
 sky130_fd_sc_hd__nor2_1 _24614_ (.A(_04705_),
    .B(_04780_),
    .Y(_04781_));
 sky130_fd_sc_hd__mux2_1 _24615_ (.A0(_04778_),
    .A1(_04781_),
    .S(_04753_),
    .X(_04782_));
 sky130_fd_sc_hd__clkbuf_1 _24616_ (.A(_04782_),
    .X(_14609_));
 sky130_fd_sc_hd__mux2_1 _24617_ (.A0(_10384_),
    .A1(_08363_),
    .S(_08472_),
    .X(_04783_));
 sky130_fd_sc_hd__clkbuf_2 _24618_ (.A(_10105_),
    .X(_04784_));
 sky130_fd_sc_hd__mux2_1 _24619_ (.A0(_04783_),
    .A1(_04769_),
    .S(_04784_),
    .X(_04785_));
 sky130_fd_sc_hd__buf_2 _24620_ (.A(_10271_),
    .X(_04786_));
 sky130_fd_sc_hd__mux4_1 _24621_ (.A0(_04785_),
    .A1(_04730_),
    .A2(_04731_),
    .A3(_04733_),
    .S0(_04786_),
    .S1(_10274_),
    .X(_04787_));
 sky130_fd_sc_hd__buf_2 _24622_ (.A(_10298_),
    .X(_04788_));
 sky130_vsdinv _24623_ (.A(_04734_),
    .Y(_04789_));
 sky130_fd_sc_hd__mux2_1 _24624_ (.A0(_04789_),
    .A1(_04738_),
    .S(_10287_),
    .X(_04790_));
 sky130_fd_sc_hd__nor2_1 _24625_ (.A(_04788_),
    .B(_04790_),
    .Y(_04791_));
 sky130_fd_sc_hd__mux2_1 _24626_ (.A0(_04787_),
    .A1(_04791_),
    .S(_04753_),
    .X(_04792_));
 sky130_fd_sc_hd__clkbuf_1 _24627_ (.A(_04792_),
    .X(_14610_));
 sky130_fd_sc_hd__mux4_1 _24628_ (.A0(_10224_),
    .A1(_10384_),
    .A2(_10214_),
    .A3(_10378_),
    .S0(_10281_),
    .S1(_04716_),
    .X(_04793_));
 sky130_fd_sc_hd__mux2_1 _24629_ (.A0(_04793_),
    .A1(_04745_),
    .S(_04701_),
    .X(_04794_));
 sky130_fd_sc_hd__mux2_1 _24630_ (.A0(_04746_),
    .A1(_04742_),
    .S(_04694_),
    .X(_04795_));
 sky130_fd_sc_hd__mux2_1 _24631_ (.A0(_04794_),
    .A1(_04795_),
    .S(_04704_),
    .X(_04796_));
 sky130_fd_sc_hd__mux2_1 _24632_ (.A0(_04743_),
    .A1(_04750_),
    .S(_04701_),
    .X(_04797_));
 sky130_fd_sc_hd__and2b_1 _24633_ (.A_N(_10274_),
    .B(_04797_),
    .X(_04798_));
 sky130_fd_sc_hd__mux2_1 _24634_ (.A0(_04796_),
    .A1(_04798_),
    .S(_04753_),
    .X(_04799_));
 sky130_fd_sc_hd__clkbuf_1 _24635_ (.A(_04799_),
    .X(_14611_));
 sky130_fd_sc_hd__mux2_1 _24636_ (.A0(_10389_),
    .A1(_10223_),
    .S(_08472_),
    .X(_04800_));
 sky130_fd_sc_hd__clkbuf_2 _24637_ (.A(_04701_),
    .X(_04801_));
 sky130_fd_sc_hd__mux4_1 _24638_ (.A0(_04800_),
    .A1(_04783_),
    .A2(_04769_),
    .A3(_04729_),
    .S0(_10285_),
    .S1(_04801_),
    .X(_04802_));
 sky130_vsdinv _24639_ (.A(_04708_),
    .Y(_04803_));
 sky130_fd_sc_hd__mux4_1 _24640_ (.A0(_04802_),
    .A1(_04702_),
    .A2(_04695_),
    .A3(_04803_),
    .S0(_04788_),
    .S1(_04755_),
    .X(_04804_));
 sky130_fd_sc_hd__clkbuf_1 _24641_ (.A(_04804_),
    .X(_14612_));
 sky130_fd_sc_hd__buf_2 _24642_ (.A(_10268_),
    .X(_04805_));
 sky130_fd_sc_hd__mux4_1 _24643_ (.A0(_10392_),
    .A1(_10389_),
    .A2(_10224_),
    .A3(_10384_),
    .S0(_04805_),
    .S1(_04764_),
    .X(_04806_));
 sky130_fd_sc_hd__buf_2 _24644_ (.A(_04722_),
    .X(_04807_));
 sky130_fd_sc_hd__mux2_1 _24645_ (.A0(_04806_),
    .A1(_04775_),
    .S(_04807_),
    .X(_04808_));
 sky130_fd_sc_hd__nor2_1 _24646_ (.A(_10273_),
    .B(_04725_),
    .Y(_04809_));
 sky130_fd_sc_hd__mux4_1 _24647_ (.A0(_04808_),
    .A1(_04720_),
    .A2(_04715_),
    .A3(_04809_),
    .S0(_04788_),
    .S1(_04755_),
    .X(_04810_));
 sky130_fd_sc_hd__clkbuf_1 _24648_ (.A(_04810_),
    .X(_14613_));
 sky130_fd_sc_hd__mux2_1 _24649_ (.A0(_10397_),
    .A1(_10392_),
    .S(_08472_),
    .X(_04811_));
 sky130_fd_sc_hd__mux2_1 _24650_ (.A0(_04811_),
    .A1(_04800_),
    .S(_04784_),
    .X(_04812_));
 sky130_fd_sc_hd__mux2_1 _24651_ (.A0(_04812_),
    .A1(_04785_),
    .S(_04807_),
    .X(_04813_));
 sky130_vsdinv _24652_ (.A(_04739_),
    .Y(_04814_));
 sky130_fd_sc_hd__buf_2 _24653_ (.A(_10275_),
    .X(_04815_));
 sky130_fd_sc_hd__clkbuf_2 _24654_ (.A(_10274_),
    .X(_04816_));
 sky130_fd_sc_hd__mux4_1 _24655_ (.A0(_04813_),
    .A1(_04735_),
    .A2(_04732_),
    .A3(_04814_),
    .S0(_04815_),
    .S1(_04816_),
    .X(_04817_));
 sky130_fd_sc_hd__clkbuf_1 _24656_ (.A(_04817_),
    .X(_14614_));
 sky130_fd_sc_hd__mux4_1 _24657_ (.A0(_10240_),
    .A1(_10397_),
    .A2(_10392_),
    .A3(_10389_),
    .S0(_04805_),
    .S1(_04764_),
    .X(_04818_));
 sky130_fd_sc_hd__mux2_1 _24658_ (.A0(_04818_),
    .A1(_04793_),
    .S(_04807_),
    .X(_04819_));
 sky130_fd_sc_hd__and2b_1 _24659_ (.A_N(_10273_),
    .B(_04750_),
    .X(_04820_));
 sky130_fd_sc_hd__mux4_1 _24660_ (.A0(_04819_),
    .A1(_04747_),
    .A2(_04744_),
    .A3(_04820_),
    .S0(_04788_),
    .S1(_04755_),
    .X(_04821_));
 sky130_fd_sc_hd__clkbuf_1 _24661_ (.A(_04821_),
    .X(_14615_));
 sky130_fd_sc_hd__mux2_1 _24662_ (.A0(_10246_),
    .A1(_10241_),
    .S(_10282_),
    .X(_04822_));
 sky130_fd_sc_hd__mux4_1 _24663_ (.A0(_04822_),
    .A1(_04811_),
    .A2(_04800_),
    .A3(_04783_),
    .S0(_10285_),
    .S1(_04801_),
    .X(_04823_));
 sky130_vsdinv _24664_ (.A(_04767_),
    .Y(_04824_));
 sky130_fd_sc_hd__mux4_1 _24665_ (.A0(_04823_),
    .A1(_04824_),
    .A2(_04771_),
    .A3(_04761_),
    .S0(_04815_),
    .S1(_04816_),
    .X(_04825_));
 sky130_fd_sc_hd__clkbuf_1 _24666_ (.A(_04825_),
    .X(_14616_));
 sky130_fd_sc_hd__mux4_1 _24667_ (.A0(_10250_),
    .A1(_10245_),
    .A2(_10240_),
    .A3(_10397_),
    .S0(_10269_),
    .S1(_04764_),
    .X(_04826_));
 sky130_fd_sc_hd__mux2_1 _24668_ (.A0(_04826_),
    .A1(_04806_),
    .S(_04757_),
    .X(_04827_));
 sky130_vsdinv _24669_ (.A(_04780_),
    .Y(_04828_));
 sky130_fd_sc_hd__mux4_1 _24670_ (.A0(_04827_),
    .A1(_04776_),
    .A2(_04777_),
    .A3(_04828_),
    .S0(_04788_),
    .S1(_04710_),
    .X(_04829_));
 sky130_fd_sc_hd__clkbuf_1 _24671_ (.A(_04829_),
    .X(_14617_));
 sky130_fd_sc_hd__mux4_1 _24672_ (.A0(_10254_),
    .A1(_10250_),
    .A2(_10246_),
    .A3(_10241_),
    .S0(_10269_),
    .S1(_10107_),
    .X(_04830_));
 sky130_fd_sc_hd__mux4_1 _24673_ (.A0(_04830_),
    .A1(_04812_),
    .A2(_04785_),
    .A3(_04730_),
    .S0(_04786_),
    .S1(_04704_),
    .X(_04831_));
 sky130_fd_sc_hd__mux2_1 _24674_ (.A0(_04731_),
    .A1(_04733_),
    .S(_10272_),
    .X(_04832_));
 sky130_fd_sc_hd__nor2_1 _24675_ (.A(_10274_),
    .B(_04832_),
    .Y(_04833_));
 sky130_fd_sc_hd__a21oi_1 _24676_ (.A1(_04788_),
    .A2(_04790_),
    .B1(_04833_),
    .Y(_04834_));
 sky130_fd_sc_hd__mux2_1 _24677_ (.A0(_04831_),
    .A1(_04834_),
    .S(_04753_),
    .X(_04835_));
 sky130_fd_sc_hd__clkbuf_1 _24678_ (.A(_04835_),
    .X(_14618_));
 sky130_fd_sc_hd__buf_2 _24679_ (.A(_10268_),
    .X(_04836_));
 sky130_fd_sc_hd__mux4_1 _24680_ (.A0(_08393_),
    .A1(_10254_),
    .A2(_08397_),
    .A3(_10245_),
    .S0(_04836_),
    .S1(_04764_),
    .X(_04837_));
 sky130_fd_sc_hd__mux2_1 _24681_ (.A0(_04837_),
    .A1(_04818_),
    .S(_04757_),
    .X(_04838_));
 sky130_fd_sc_hd__buf_2 _24682_ (.A(_04762_),
    .X(_04839_));
 sky130_fd_sc_hd__mux4_1 _24683_ (.A0(_04838_),
    .A1(_04795_),
    .A2(_04794_),
    .A3(_04797_),
    .S0(_04815_),
    .S1(_04839_),
    .X(_04840_));
 sky130_fd_sc_hd__clkbuf_1 _24684_ (.A(_04840_),
    .X(_14619_));
 sky130_fd_sc_hd__o21ai_1 _24685_ (.A1(_08757_),
    .A2(_08470_),
    .B1(_04707_),
    .Y(_04841_));
 sky130_fd_sc_hd__mux2_1 _24686_ (.A0(_10331_),
    .A1(_10334_),
    .S(_10282_),
    .X(_04842_));
 sky130_fd_sc_hd__mux2_1 _24687_ (.A0(_10311_),
    .A1(_10322_),
    .S(_10282_),
    .X(_04843_));
 sky130_fd_sc_hd__mux2_1 _24688_ (.A0(_10337_),
    .A1(_08461_),
    .S(_10269_),
    .X(_04844_));
 sky130_fd_sc_hd__mux4_1 _24689_ (.A0(_04841_),
    .A1(_04842_),
    .A2(_04843_),
    .A3(_04844_),
    .S0(_04706_),
    .S1(_10108_),
    .X(_04845_));
 sky130_fd_sc_hd__mux2_1 _24690_ (.A0(_10367_),
    .A1(_10197_),
    .S(_04805_),
    .X(_04846_));
 sky130_fd_sc_hd__mux2_1 _24691_ (.A0(_10372_),
    .A1(_10206_),
    .S(_04805_),
    .X(_04847_));
 sky130_fd_sc_hd__mux2_1 _24692_ (.A0(_08355_),
    .A1(_08363_),
    .S(_04749_),
    .X(_04848_));
 sky130_fd_sc_hd__mux2_1 _24693_ (.A0(_08359_),
    .A1(_10223_),
    .S(_10281_),
    .X(_04849_));
 sky130_fd_sc_hd__clkbuf_4 _24694_ (.A(_10106_),
    .X(_04850_));
 sky130_fd_sc_hd__mux4_2 _24695_ (.A0(_04846_),
    .A1(_04847_),
    .A2(_04848_),
    .A3(_04849_),
    .S0(_04850_),
    .S1(_04757_),
    .X(_04851_));
 sky130_fd_sc_hd__mux2_1 _24696_ (.A0(_10344_),
    .A1(_10157_),
    .S(_04836_),
    .X(_04852_));
 sky130_fd_sc_hd__mux2_1 _24697_ (.A0(_10163_),
    .A1(_08412_),
    .S(_04836_),
    .X(_04853_));
 sky130_fd_sc_hd__mux2_1 _24698_ (.A0(_10354_),
    .A1(_10357_),
    .S(_04805_),
    .X(_04854_));
 sky130_fd_sc_hd__mux2_1 _24699_ (.A0(_10361_),
    .A1(_10187_),
    .S(_04836_),
    .X(_04855_));
 sky130_fd_sc_hd__mux4_1 _24700_ (.A0(_04852_),
    .A1(_04853_),
    .A2(_04854_),
    .A3(_04855_),
    .S0(_04758_),
    .S1(_04807_),
    .X(_04856_));
 sky130_fd_sc_hd__mux2_1 _24701_ (.A0(_08423_),
    .A1(_10232_),
    .S(_04718_),
    .X(_04857_));
 sky130_fd_sc_hd__mux2_1 _24702_ (.A0(_10396_),
    .A1(_10240_),
    .S(_10281_),
    .X(_04858_));
 sky130_fd_sc_hd__mux2_1 _24703_ (.A0(_04857_),
    .A1(_04858_),
    .S(_10284_),
    .X(_04859_));
 sky130_fd_sc_hd__mux2_1 _24704_ (.A0(_10245_),
    .A1(_08397_),
    .S(_04718_),
    .X(_04860_));
 sky130_fd_sc_hd__mux2_1 _24705_ (.A0(_10254_),
    .A1(net291),
    .S(_04718_),
    .X(_04861_));
 sky130_fd_sc_hd__mux2_1 _24706_ (.A0(_04860_),
    .A1(_04861_),
    .S(_10284_),
    .X(_04862_));
 sky130_fd_sc_hd__mux2_2 _24707_ (.A0(_04859_),
    .A1(_04862_),
    .S(_04786_),
    .X(_04863_));
 sky130_fd_sc_hd__mux4_1 _24708_ (.A0(_04845_),
    .A1(_04851_),
    .A2(_04856_),
    .A3(_04863_),
    .S0(_04815_),
    .S1(_04839_),
    .X(_04864_));
 sky130_fd_sc_hd__clkbuf_1 _24709_ (.A(_04864_),
    .X(_14620_));
 sky130_fd_sc_hd__mux2_1 _24710_ (.A0(_10104_),
    .A1(_10311_),
    .S(_10282_),
    .X(_04865_));
 sky130_fd_sc_hd__mux2_1 _24711_ (.A0(_10334_),
    .A1(_10337_),
    .S(_10269_),
    .X(_04866_));
 sky130_fd_sc_hd__mux2_1 _24712_ (.A0(_10322_),
    .A1(_10331_),
    .S(_10282_),
    .X(_04867_));
 sky130_fd_sc_hd__mux2_1 _24713_ (.A0(_08461_),
    .A1(_10344_),
    .S(_10269_),
    .X(_04868_));
 sky130_fd_sc_hd__clkbuf_2 _24714_ (.A(_10107_),
    .X(_04869_));
 sky130_fd_sc_hd__mux4_1 _24715_ (.A0(_04865_),
    .A1(_04866_),
    .A2(_04867_),
    .A3(_04868_),
    .S0(_04706_),
    .S1(_04869_),
    .X(_04870_));
 sky130_fd_sc_hd__mux2_1 _24716_ (.A0(_08382_),
    .A1(_08351_),
    .S(_08472_),
    .X(_04871_));
 sky130_fd_sc_hd__mux2_1 _24717_ (.A0(_08374_),
    .A1(_08355_),
    .S(_04749_),
    .X(_04872_));
 sky130_fd_sc_hd__mux2_1 _24718_ (.A0(_08363_),
    .A1(_08359_),
    .S(_04749_),
    .X(_04873_));
 sky130_fd_sc_hd__mux2_1 _24719_ (.A0(_10223_),
    .A1(_08423_),
    .S(_04696_),
    .X(_04874_));
 sky130_fd_sc_hd__mux4_2 _24720_ (.A0(_04871_),
    .A1(_04872_),
    .A2(_04873_),
    .A3(_04874_),
    .S0(_04850_),
    .S1(_04757_),
    .X(_04875_));
 sky130_fd_sc_hd__mux2_1 _24721_ (.A0(_10157_),
    .A1(_10163_),
    .S(_04836_),
    .X(_04876_));
 sky130_fd_sc_hd__mux2_1 _24722_ (.A0(_08412_),
    .A1(_10354_),
    .S(_04805_),
    .X(_04877_));
 sky130_fd_sc_hd__mux2_1 _24723_ (.A0(_10357_),
    .A1(_10361_),
    .S(_04836_),
    .X(_04878_));
 sky130_fd_sc_hd__mux2_1 _24724_ (.A0(_10187_),
    .A1(_10367_),
    .S(_08472_),
    .X(_04879_));
 sky130_fd_sc_hd__mux4_1 _24725_ (.A0(_04876_),
    .A1(_04877_),
    .A2(_04878_),
    .A3(_04879_),
    .S0(_04758_),
    .S1(_04807_),
    .X(_04880_));
 sky130_fd_sc_hd__mux2_1 _24726_ (.A0(_10232_),
    .A1(_10396_),
    .S(_04696_),
    .X(_04881_));
 sky130_fd_sc_hd__mux2_1 _24727_ (.A0(_10240_),
    .A1(_10245_),
    .S(_04696_),
    .X(_04882_));
 sky130_fd_sc_hd__mux2_1 _24728_ (.A0(_04881_),
    .A1(_04882_),
    .S(_10284_),
    .X(_04883_));
 sky130_fd_sc_hd__mux2_1 _24729_ (.A0(net288),
    .A1(_10254_),
    .S(_04686_),
    .X(_04884_));
 sky130_fd_sc_hd__o21ai_4 _24730_ (.A1(instr_sra),
    .A2(instr_srai),
    .B1(net291),
    .Y(_04885_));
 sky130_fd_sc_hd__nand2_1 _24731_ (.A(_10106_),
    .B(_04885_),
    .Y(_04886_));
 sky130_fd_sc_hd__and2_1 _24732_ (.A(net291),
    .B(_08470_),
    .X(_04887_));
 sky130_fd_sc_hd__o22a_1 _24733_ (.A1(_04764_),
    .A2(_04884_),
    .B1(_04886_),
    .B2(_04887_),
    .X(_04888_));
 sky130_fd_sc_hd__mux2_2 _24734_ (.A0(_04883_),
    .A1(_04888_),
    .S(_04786_),
    .X(_04889_));
 sky130_fd_sc_hd__mux4_1 _24735_ (.A0(_04870_),
    .A1(_04875_),
    .A2(_04880_),
    .A3(_04889_),
    .S0(_04815_),
    .S1(_04839_),
    .X(_04890_));
 sky130_fd_sc_hd__clkbuf_1 _24736_ (.A(_04890_),
    .X(_14631_));
 sky130_fd_sc_hd__mux4_1 _24737_ (.A0(_04843_),
    .A1(_04844_),
    .A2(_04842_),
    .A3(_04852_),
    .S0(_04706_),
    .S1(_04869_),
    .X(_04891_));
 sky130_fd_sc_hd__mux4_1 _24738_ (.A0(_04853_),
    .A1(_04854_),
    .A2(_04855_),
    .A3(_04846_),
    .S0(_04850_),
    .S1(_04757_),
    .X(_04892_));
 sky130_fd_sc_hd__mux4_2 _24739_ (.A0(_04847_),
    .A1(_04848_),
    .A2(_04849_),
    .A3(_04857_),
    .S0(_04850_),
    .S1(_04770_),
    .X(_04893_));
 sky130_fd_sc_hd__mux2_1 _24740_ (.A0(_04858_),
    .A1(_04860_),
    .S(_04784_),
    .X(_04894_));
 sky130_fd_sc_hd__o21a_1 _24741_ (.A1(_10107_),
    .A2(_04861_),
    .B1(_04886_),
    .X(_04895_));
 sky130_fd_sc_hd__mux2_2 _24742_ (.A0(_04894_),
    .A1(_04895_),
    .S(_04786_),
    .X(_04896_));
 sky130_fd_sc_hd__mux4_1 _24743_ (.A0(_04891_),
    .A1(_04892_),
    .A2(_04893_),
    .A3(_04896_),
    .S0(_04762_),
    .S1(_04710_),
    .X(_04897_));
 sky130_fd_sc_hd__clkbuf_1 _24744_ (.A(_04897_),
    .X(_14642_));
 sky130_fd_sc_hd__mux4_1 _24745_ (.A0(_04867_),
    .A1(_04868_),
    .A2(_04866_),
    .A3(_04876_),
    .S0(_04706_),
    .S1(_04869_),
    .X(_04898_));
 sky130_fd_sc_hd__mux4_2 _24746_ (.A0(_04872_),
    .A1(_04873_),
    .A2(_04874_),
    .A3(_04881_),
    .S0(_04850_),
    .S1(_04770_),
    .X(_04899_));
 sky130_fd_sc_hd__mux4_1 _24747_ (.A0(_04877_),
    .A1(_04878_),
    .A2(_04879_),
    .A3(_04871_),
    .S0(_04850_),
    .S1(_04807_),
    .X(_04900_));
 sky130_fd_sc_hd__mux2_1 _24748_ (.A0(_04882_),
    .A1(_04884_),
    .S(_04692_),
    .X(_04901_));
 sky130_fd_sc_hd__o21a_1 _24749_ (.A1(instr_sra),
    .A2(instr_srai),
    .B1(_08393_),
    .X(_04902_));
 sky130_fd_sc_hd__o21a_1 _24750_ (.A1(_04887_),
    .A2(_04902_),
    .B1(_04886_),
    .X(_04903_));
 sky130_fd_sc_hd__mux2_2 _24751_ (.A0(_04901_),
    .A1(_04903_),
    .S(_04786_),
    .X(_04904_));
 sky130_fd_sc_hd__buf_2 _24752_ (.A(_10275_),
    .X(_04905_));
 sky130_fd_sc_hd__mux4_1 _24753_ (.A0(_04898_),
    .A1(_04899_),
    .A2(_04900_),
    .A3(_04904_),
    .S0(_04905_),
    .S1(_04839_),
    .X(_04906_));
 sky130_fd_sc_hd__clkbuf_1 _24754_ (.A(_04906_),
    .X(_14645_));
 sky130_fd_sc_hd__mux4_1 _24755_ (.A0(_04842_),
    .A1(_04844_),
    .A2(_04852_),
    .A3(_04853_),
    .S0(_10285_),
    .S1(_04801_),
    .X(_04907_));
 sky130_fd_sc_hd__mux2_1 _24756_ (.A0(_04848_),
    .A1(_04849_),
    .S(_04784_),
    .X(_04908_));
 sky130_fd_sc_hd__mux2_1 _24757_ (.A0(_04908_),
    .A1(_04859_),
    .S(_04770_),
    .X(_04909_));
 sky130_fd_sc_hd__mux4_1 _24758_ (.A0(_04854_),
    .A1(_04846_),
    .A2(_04855_),
    .A3(_04847_),
    .S0(_10272_),
    .S1(_04869_),
    .X(_04910_));
 sky130_fd_sc_hd__nand2_1 _24759_ (.A(_10287_),
    .B(_04885_),
    .Y(_04911_));
 sky130_fd_sc_hd__o21a_1 _24760_ (.A1(_04723_),
    .A2(_04862_),
    .B1(_04911_),
    .X(_04912_));
 sky130_fd_sc_hd__mux4_1 _24761_ (.A0(_04907_),
    .A1(_04909_),
    .A2(_04910_),
    .A3(_04912_),
    .S0(_04905_),
    .S1(_04839_),
    .X(_04913_));
 sky130_fd_sc_hd__clkbuf_1 _24762_ (.A(_04913_),
    .X(_14646_));
 sky130_fd_sc_hd__mux4_1 _24763_ (.A0(_04866_),
    .A1(_04868_),
    .A2(_04876_),
    .A3(_04877_),
    .S0(_04758_),
    .S1(_04801_),
    .X(_04914_));
 sky130_fd_sc_hd__mux2_1 _24764_ (.A0(_04873_),
    .A1(_04874_),
    .S(_04784_),
    .X(_04915_));
 sky130_fd_sc_hd__mux2_1 _24765_ (.A0(_04915_),
    .A1(_04883_),
    .S(_04770_),
    .X(_04916_));
 sky130_fd_sc_hd__mux4_1 _24766_ (.A0(_04878_),
    .A1(_04871_),
    .A2(_04879_),
    .A3(_04872_),
    .S0(_10272_),
    .S1(_04869_),
    .X(_04917_));
 sky130_fd_sc_hd__o21a_1 _24767_ (.A1(_04723_),
    .A2(_04888_),
    .B1(_04911_),
    .X(_04918_));
 sky130_fd_sc_hd__mux4_1 _24768_ (.A0(_04914_),
    .A1(_04916_),
    .A2(_04917_),
    .A3(_04918_),
    .S0(_04905_),
    .S1(_04839_),
    .X(_04919_));
 sky130_fd_sc_hd__clkbuf_1 _24769_ (.A(_04919_),
    .X(_14647_));
 sky130_fd_sc_hd__mux4_1 _24770_ (.A0(_04844_),
    .A1(_04852_),
    .A2(_04853_),
    .A3(_04854_),
    .S0(_04758_),
    .S1(_04801_),
    .X(_04920_));
 sky130_fd_sc_hd__mux2_1 _24771_ (.A0(_04849_),
    .A1(_04857_),
    .S(_04784_),
    .X(_04921_));
 sky130_fd_sc_hd__mux2_1 _24772_ (.A0(_04921_),
    .A1(_04894_),
    .S(_04770_),
    .X(_04922_));
 sky130_fd_sc_hd__mux4_1 _24773_ (.A0(_04855_),
    .A1(_04847_),
    .A2(_04846_),
    .A3(_04848_),
    .S0(_10272_),
    .S1(_04869_),
    .X(_04923_));
 sky130_fd_sc_hd__o21a_1 _24774_ (.A1(_04723_),
    .A2(_04895_),
    .B1(_04911_),
    .X(_04924_));
 sky130_fd_sc_hd__clkbuf_2 _24775_ (.A(_04762_),
    .X(_04925_));
 sky130_fd_sc_hd__mux4_1 _24776_ (.A0(_04920_),
    .A1(_04922_),
    .A2(_04923_),
    .A3(_04924_),
    .S0(_04905_),
    .S1(_04925_),
    .X(_04926_));
 sky130_fd_sc_hd__clkbuf_1 _24777_ (.A(_04926_),
    .X(_14648_));
 sky130_fd_sc_hd__mux4_1 _24778_ (.A0(_04868_),
    .A1(_04876_),
    .A2(_04877_),
    .A3(_04878_),
    .S0(_04758_),
    .S1(_04801_),
    .X(_04927_));
 sky130_fd_sc_hd__mux2_1 _24779_ (.A0(_04874_),
    .A1(_04881_),
    .S(_04712_),
    .X(_04928_));
 sky130_fd_sc_hd__mux2_1 _24780_ (.A0(_04928_),
    .A1(_04901_),
    .S(_04694_),
    .X(_04929_));
 sky130_fd_sc_hd__mux4_1 _24781_ (.A0(_04879_),
    .A1(_04872_),
    .A2(_04871_),
    .A3(_04873_),
    .S0(_10271_),
    .S1(_10107_),
    .X(_04930_));
 sky130_fd_sc_hd__and2_1 _24782_ (.A(_04903_),
    .B(_04911_),
    .X(_04931_));
 sky130_fd_sc_hd__mux4_1 _24783_ (.A0(_04927_),
    .A1(_04929_),
    .A2(_04930_),
    .A3(_04931_),
    .S0(_04905_),
    .S1(_04925_),
    .X(_04932_));
 sky130_fd_sc_hd__clkbuf_1 _24784_ (.A(_04932_),
    .X(_14649_));
 sky130_fd_sc_hd__buf_1 _24785_ (.A(_04902_),
    .X(_04933_));
 sky130_fd_sc_hd__mux4_1 _24786_ (.A0(_04856_),
    .A1(_04863_),
    .A2(_04851_),
    .A3(_04933_),
    .S0(_04905_),
    .S1(_04925_),
    .X(_04934_));
 sky130_fd_sc_hd__clkbuf_1 _24787_ (.A(_04934_),
    .X(_14650_));
 sky130_fd_sc_hd__buf_2 _24788_ (.A(_10275_),
    .X(_04935_));
 sky130_fd_sc_hd__mux4_1 _24789_ (.A0(_04880_),
    .A1(_04889_),
    .A2(_04875_),
    .A3(_04933_),
    .S0(_04935_),
    .S1(_04925_),
    .X(_04936_));
 sky130_fd_sc_hd__clkbuf_1 _24790_ (.A(_04936_),
    .X(_14651_));
 sky130_fd_sc_hd__mux4_1 _24791_ (.A0(_04892_),
    .A1(_04893_),
    .A2(_04896_),
    .A3(_04933_),
    .S0(_04762_),
    .S1(_04710_),
    .X(_04937_));
 sky130_fd_sc_hd__clkbuf_1 _24792_ (.A(_04937_),
    .X(_14621_));
 sky130_fd_sc_hd__mux4_1 _24793_ (.A0(_04900_),
    .A1(_04904_),
    .A2(_04899_),
    .A3(_04933_),
    .S0(_04935_),
    .S1(_04925_),
    .X(_04938_));
 sky130_fd_sc_hd__clkbuf_1 _24794_ (.A(_04938_),
    .X(_14622_));
 sky130_fd_sc_hd__mux4_1 _24795_ (.A0(_04910_),
    .A1(_04912_),
    .A2(_04909_),
    .A3(_04933_),
    .S0(_04935_),
    .S1(_04925_),
    .X(_04939_));
 sky130_fd_sc_hd__clkbuf_1 _24796_ (.A(_04939_),
    .X(_14623_));
 sky130_fd_sc_hd__mux4_1 _24797_ (.A0(_04917_),
    .A1(_04918_),
    .A2(_04916_),
    .A3(_04933_),
    .S0(_04935_),
    .S1(_04768_),
    .X(_04940_));
 sky130_fd_sc_hd__clkbuf_1 _24798_ (.A(_04940_),
    .X(_14624_));
 sky130_fd_sc_hd__mux4_1 _24799_ (.A0(_04923_),
    .A1(_04924_),
    .A2(_04922_),
    .A3(_04902_),
    .S0(_04935_),
    .S1(_04768_),
    .X(_04941_));
 sky130_fd_sc_hd__clkbuf_1 _24800_ (.A(_04941_),
    .X(_14625_));
 sky130_fd_sc_hd__mux2_1 _24801_ (.A0(_04930_),
    .A1(_04929_),
    .S(_04704_),
    .X(_04942_));
 sky130_fd_sc_hd__nand2_1 _24802_ (.A(_10298_),
    .B(_04885_),
    .Y(_04943_));
 sky130_fd_sc_hd__and3_1 _24803_ (.A(_04903_),
    .B(_04911_),
    .C(_04943_),
    .X(_04944_));
 sky130_fd_sc_hd__mux2_1 _24804_ (.A0(_04942_),
    .A1(_04944_),
    .S(_04753_),
    .X(_04945_));
 sky130_fd_sc_hd__clkbuf_1 _24805_ (.A(_04945_),
    .X(_14626_));
 sky130_fd_sc_hd__clkbuf_2 _24806_ (.A(_10276_),
    .X(_04946_));
 sky130_fd_sc_hd__clkbuf_2 _24807_ (.A(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__mux2_1 _24808_ (.A0(_04851_),
    .A1(_04863_),
    .S(_04768_),
    .X(_04948_));
 sky130_fd_sc_hd__nand2_2 _24809_ (.A(_04935_),
    .B(_04885_),
    .Y(_04949_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _24810_ (.A(_04949_),
    .X(_04950_));
 sky130_fd_sc_hd__o21a_1 _24811_ (.A1(_04947_),
    .A2(_04948_),
    .B1(_04950_),
    .X(_14627_));
 sky130_fd_sc_hd__mux2_1 _24812_ (.A0(_04875_),
    .A1(_04889_),
    .S(_04768_),
    .X(_04951_));
 sky130_fd_sc_hd__o21a_1 _24813_ (.A1(_04947_),
    .A2(_04951_),
    .B1(_04950_),
    .X(_14628_));
 sky130_fd_sc_hd__clkbuf_2 _24814_ (.A(_10298_),
    .X(_04952_));
 sky130_fd_sc_hd__mux2_1 _24815_ (.A0(_04893_),
    .A1(_04896_),
    .S(_04952_),
    .X(_04953_));
 sky130_fd_sc_hd__o21a_1 _24816_ (.A1(_04947_),
    .A2(_04953_),
    .B1(_04950_),
    .X(_14629_));
 sky130_fd_sc_hd__mux2_1 _24817_ (.A0(_04899_),
    .A1(_04904_),
    .S(_04952_),
    .X(_04954_));
 sky130_fd_sc_hd__o21a_1 _24818_ (.A1(_04947_),
    .A2(_04954_),
    .B1(_04950_),
    .X(_14630_));
 sky130_fd_sc_hd__mux2_1 _24819_ (.A0(_04909_),
    .A1(_04912_),
    .S(_04952_),
    .X(_04955_));
 sky130_fd_sc_hd__o21a_1 _24820_ (.A1(_04947_),
    .A2(_04955_),
    .B1(_04950_),
    .X(_14632_));
 sky130_fd_sc_hd__mux2_1 _24821_ (.A0(_04916_),
    .A1(_04918_),
    .S(_04952_),
    .X(_04956_));
 sky130_fd_sc_hd__o21a_1 _24822_ (.A1(_04947_),
    .A2(_04956_),
    .B1(_04950_),
    .X(_14633_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _24823_ (.A(_04946_),
    .X(_04957_));
 sky130_fd_sc_hd__mux2_1 _24824_ (.A0(_04922_),
    .A1(_04924_),
    .S(_04952_),
    .X(_04958_));
 sky130_fd_sc_hd__clkbuf_2 _24825_ (.A(_04949_),
    .X(_04959_));
 sky130_fd_sc_hd__o21a_1 _24826_ (.A1(_04957_),
    .A2(_04958_),
    .B1(_04959_),
    .X(_14634_));
 sky130_fd_sc_hd__mux2_1 _24827_ (.A0(_04929_),
    .A1(_04931_),
    .S(_04952_),
    .X(_04960_));
 sky130_fd_sc_hd__o21a_1 _24828_ (.A1(_04957_),
    .A2(_04960_),
    .B1(_04959_),
    .X(_14635_));
 sky130_fd_sc_hd__buf_4 _24829_ (.A(_04762_),
    .X(_04961_));
 sky130_fd_sc_hd__clkbuf_2 _24830_ (.A(_04943_),
    .X(_04962_));
 sky130_fd_sc_hd__o21a_1 _24831_ (.A1(_04961_),
    .A2(_04863_),
    .B1(_04962_),
    .X(_04963_));
 sky130_fd_sc_hd__o21a_1 _24832_ (.A1(_04957_),
    .A2(_04963_),
    .B1(_04959_),
    .X(_14636_));
 sky130_fd_sc_hd__o21a_1 _24833_ (.A1(_04961_),
    .A2(_04889_),
    .B1(_04962_),
    .X(_04964_));
 sky130_fd_sc_hd__o21a_1 _24834_ (.A1(_04957_),
    .A2(_04964_),
    .B1(_04959_),
    .X(_14637_));
 sky130_fd_sc_hd__o21a_1 _24835_ (.A1(_04961_),
    .A2(_04896_),
    .B1(_04962_),
    .X(_04965_));
 sky130_fd_sc_hd__o21a_1 _24836_ (.A1(_04957_),
    .A2(_04965_),
    .B1(_04959_),
    .X(_14638_));
 sky130_fd_sc_hd__o21a_1 _24837_ (.A1(_04816_),
    .A2(_04904_),
    .B1(_04962_),
    .X(_04966_));
 sky130_fd_sc_hd__o21a_1 _24838_ (.A1(_04957_),
    .A2(_04966_),
    .B1(_04959_),
    .X(_14639_));
 sky130_fd_sc_hd__o21a_1 _24839_ (.A1(_04816_),
    .A2(_04912_),
    .B1(_04962_),
    .X(_04967_));
 sky130_fd_sc_hd__o21a_1 _24840_ (.A1(_04756_),
    .A2(_04967_),
    .B1(_04949_),
    .X(_14640_));
 sky130_fd_sc_hd__o21a_1 _24841_ (.A1(_04816_),
    .A2(_04918_),
    .B1(_04962_),
    .X(_04968_));
 sky130_fd_sc_hd__o21a_1 _24842_ (.A1(_04756_),
    .A2(_04968_),
    .B1(_04949_),
    .X(_14641_));
 sky130_fd_sc_hd__o21a_1 _24843_ (.A1(_04816_),
    .A2(_04924_),
    .B1(_04943_),
    .X(_04969_));
 sky130_fd_sc_hd__o21a_1 _24844_ (.A1(_04756_),
    .A2(_04969_),
    .B1(_04949_),
    .X(_14643_));
 sky130_fd_sc_hd__and2_1 _24845_ (.A(_04944_),
    .B(_04949_),
    .X(_04970_));
 sky130_fd_sc_hd__clkbuf_1 _24846_ (.A(_04970_),
    .X(_14644_));
 sky130_fd_sc_hd__clkbuf_2 _24847_ (.A(\irq_state[0] ),
    .X(_04971_));
 sky130_fd_sc_hd__clkbuf_2 _24848_ (.A(_04971_),
    .X(_04972_));
 sky130_fd_sc_hd__and2b_1 _24849_ (.A_N(_10316_),
    .B(_10317_),
    .X(_04973_));
 sky130_fd_sc_hd__nor2_2 _24850_ (.A(_08278_),
    .B(_04973_),
    .Y(_04974_));
 sky130_fd_sc_hd__clkbuf_2 _24851_ (.A(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__o21a_1 _24852_ (.A1(_04972_),
    .A2(_04975_),
    .B1(\reg_next_pc[0] ),
    .X(_04976_));
 sky130_fd_sc_hd__buf_2 _24853_ (.A(_10304_),
    .X(_04977_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _24854_ (.A(_04973_),
    .X(_04978_));
 sky130_fd_sc_hd__clkbuf_2 _24855_ (.A(latched_stalu),
    .X(_04979_));
 sky130_fd_sc_hd__clkbuf_2 _24856_ (.A(_04979_),
    .X(_04980_));
 sky130_fd_sc_hd__buf_2 _24857_ (.A(_04980_),
    .X(_04981_));
 sky130_fd_sc_hd__clkbuf_2 _24858_ (.A(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__clkbuf_2 _24859_ (.A(_04982_),
    .X(_04983_));
 sky130_fd_sc_hd__buf_2 _24860_ (.A(_04983_),
    .X(_04984_));
 sky130_fd_sc_hd__mux2_1 _24861_ (.A0(\reg_out[0] ),
    .A1(\alu_out_q[0] ),
    .S(_04984_),
    .X(_04985_));
 sky130_fd_sc_hd__a22o_1 _24862_ (.A1(_04977_),
    .A2(_08240_),
    .B1(_04978_),
    .B2(_04985_),
    .X(_04986_));
 sky130_fd_sc_hd__or2_4 _24863_ (.A(_04976_),
    .B(_04986_),
    .X(_04987_));
 sky130_fd_sc_hd__clkbuf_2 _24864_ (.A(_04987_),
    .X(_04988_));
 sky130_fd_sc_hd__o31ai_4 _24865_ (.A1(_10316_),
    .A2(_10317_),
    .A3(_08278_),
    .B1(_08175_),
    .Y(_04989_));
 sky130_fd_sc_hd__or3_2 _24866_ (.A(\latched_rd[1] ),
    .B(\latched_rd[0] ),
    .C(_04989_),
    .X(_04990_));
 sky130_fd_sc_hd__or3b_2 _24867_ (.A(\latched_rd[4] ),
    .B(\latched_rd[3] ),
    .C_N(\latched_rd[2] ),
    .X(_04991_));
 sky130_fd_sc_hd__nor2_1 _24868_ (.A(_04990_),
    .B(_04991_),
    .Y(_04992_));
 sky130_fd_sc_hd__clkbuf_4 _24869_ (.A(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__buf_2 _24870_ (.A(_04993_),
    .X(_04994_));
 sky130_fd_sc_hd__mux2_1 _24871_ (.A0(\cpuregs[4][0] ),
    .A1(_04988_),
    .S(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__clkbuf_1 _24872_ (.A(_04995_),
    .X(_00114_));
 sky130_fd_sc_hd__or2_1 _24873_ (.A(_08278_),
    .B(_04973_),
    .X(_04996_));
 sky130_fd_sc_hd__buf_2 _24874_ (.A(_04996_),
    .X(_04997_));
 sky130_fd_sc_hd__clkbuf_2 _24875_ (.A(_04973_),
    .X(_04998_));
 sky130_fd_sc_hd__clkbuf_2 _24876_ (.A(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__mux2_1 _24877_ (.A0(\reg_out[1] ),
    .A1(\alu_out_q[1] ),
    .S(_04979_),
    .X(_05000_));
 sky130_fd_sc_hd__and2_1 _24878_ (.A(_04999_),
    .B(_05000_),
    .X(_05001_));
 sky130_fd_sc_hd__clkbuf_2 _24879_ (.A(_04971_),
    .X(_05002_));
 sky130_fd_sc_hd__clkbuf_2 _24880_ (.A(_10304_),
    .X(_05003_));
 sky130_fd_sc_hd__a221o_1 _24881_ (.A1(_05002_),
    .A2(\reg_next_pc[1] ),
    .B1(_08263_),
    .B2(_05003_),
    .C1(_04975_),
    .X(_05004_));
 sky130_fd_sc_hd__o22a_2 _24882_ (.A1(_08184_),
    .A2(_04997_),
    .B1(_05001_),
    .B2(_05004_),
    .X(_05005_));
 sky130_fd_sc_hd__clkbuf_2 _24883_ (.A(_05005_),
    .X(_05006_));
 sky130_fd_sc_hd__mux2_1 _24884_ (.A0(\cpuregs[4][1] ),
    .A1(_05006_),
    .S(_04994_),
    .X(_05007_));
 sky130_fd_sc_hd__clkbuf_1 _24885_ (.A(_05007_),
    .X(_00115_));
 sky130_fd_sc_hd__buf_2 _24886_ (.A(\reg_pc[2] ),
    .X(_05008_));
 sky130_fd_sc_hd__clkbuf_4 _24887_ (.A(_04974_),
    .X(_05009_));
 sky130_fd_sc_hd__mux2_1 _24888_ (.A0(\reg_out[2] ),
    .A1(\alu_out_q[2] ),
    .S(latched_stalu),
    .X(_05010_));
 sky130_fd_sc_hd__clkbuf_2 _24889_ (.A(_10304_),
    .X(_05011_));
 sky130_fd_sc_hd__clkbuf_2 _24890_ (.A(_04974_),
    .X(_05012_));
 sky130_fd_sc_hd__a221o_1 _24891_ (.A1(_05002_),
    .A2(\reg_next_pc[2] ),
    .B1(_08268_),
    .B2(_05011_),
    .C1(_05012_),
    .X(_05013_));
 sky130_fd_sc_hd__a21oi_1 _24892_ (.A1(_04999_),
    .A2(_05010_),
    .B1(_05013_),
    .Y(_05014_));
 sky130_fd_sc_hd__a21oi_4 _24893_ (.A1(_05008_),
    .A2(_05009_),
    .B1(_05014_),
    .Y(_05015_));
 sky130_fd_sc_hd__clkbuf_2 _24894_ (.A(_05015_),
    .X(_05016_));
 sky130_fd_sc_hd__mux2_1 _24895_ (.A0(\cpuregs[4][2] ),
    .A1(_05016_),
    .S(_04994_),
    .X(_05017_));
 sky130_fd_sc_hd__clkbuf_1 _24896_ (.A(_05017_),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _24897_ (.A0(\reg_out[3] ),
    .A1(\alu_out_q[3] ),
    .S(latched_stalu),
    .X(_05018_));
 sky130_fd_sc_hd__and2_1 _24898_ (.A(_04978_),
    .B(_05018_),
    .X(_05019_));
 sky130_fd_sc_hd__a221o_1 _24899_ (.A1(_05002_),
    .A2(\reg_next_pc[3] ),
    .B1(_08236_),
    .B2(_05003_),
    .C1(_04975_),
    .X(_05020_));
 sky130_fd_sc_hd__xor2_1 _24900_ (.A(_08874_),
    .B(_05008_),
    .X(_05021_));
 sky130_fd_sc_hd__o22a_2 _24901_ (.A1(_05019_),
    .A2(_05020_),
    .B1(_05021_),
    .B2(_04997_),
    .X(_05022_));
 sky130_fd_sc_hd__clkbuf_2 _24902_ (.A(_05022_),
    .X(_05023_));
 sky130_fd_sc_hd__mux2_1 _24903_ (.A0(\cpuregs[4][3] ),
    .A1(_05023_),
    .S(_04994_),
    .X(_05024_));
 sky130_fd_sc_hd__clkbuf_1 _24904_ (.A(_05024_),
    .X(_00117_));
 sky130_fd_sc_hd__and2_1 _24905_ (.A(_04972_),
    .B(\reg_next_pc[4] ),
    .X(_05025_));
 sky130_fd_sc_hd__mux2_1 _24906_ (.A0(\reg_out[4] ),
    .A1(\alu_out_q[4] ),
    .S(_04979_),
    .X(_05026_));
 sky130_fd_sc_hd__a221o_1 _24907_ (.A1(_05003_),
    .A2(_08267_),
    .B1(_04978_),
    .B2(_05026_),
    .C1(_04975_),
    .X(_05027_));
 sky130_fd_sc_hd__and3_1 _24908_ (.A(\reg_pc[4] ),
    .B(_08874_),
    .C(_05008_),
    .X(_05028_));
 sky130_fd_sc_hd__a21oi_1 _24909_ (.A1(_08874_),
    .A2(_05008_),
    .B1(\reg_pc[4] ),
    .Y(_05029_));
 sky130_fd_sc_hd__nor2_1 _24910_ (.A(_05028_),
    .B(_05029_),
    .Y(_05030_));
 sky130_fd_sc_hd__o22a_2 _24911_ (.A1(_05025_),
    .A2(_05027_),
    .B1(_05030_),
    .B2(_04997_),
    .X(_05031_));
 sky130_fd_sc_hd__clkbuf_2 _24912_ (.A(_05031_),
    .X(_05032_));
 sky130_fd_sc_hd__mux2_1 _24913_ (.A0(\cpuregs[4][4] ),
    .A1(_05032_),
    .S(_04994_),
    .X(_05033_));
 sky130_fd_sc_hd__clkbuf_1 _24914_ (.A(_05033_),
    .X(_00118_));
 sky130_fd_sc_hd__mux2_1 _24915_ (.A0(\reg_out[5] ),
    .A1(\alu_out_q[5] ),
    .S(_04979_),
    .X(_05034_));
 sky130_fd_sc_hd__and2_1 _24916_ (.A(_04978_),
    .B(_05034_),
    .X(_05035_));
 sky130_fd_sc_hd__a221o_1 _24917_ (.A1(_05002_),
    .A2(\reg_next_pc[5] ),
    .B1(_08265_),
    .B2(_05003_),
    .C1(_04975_),
    .X(_05036_));
 sky130_fd_sc_hd__and2_1 _24918_ (.A(\reg_pc[5] ),
    .B(_05028_),
    .X(_05037_));
 sky130_fd_sc_hd__nor2_1 _24919_ (.A(\reg_pc[5] ),
    .B(_05028_),
    .Y(_05038_));
 sky130_fd_sc_hd__nor2_1 _24920_ (.A(_05037_),
    .B(_05038_),
    .Y(_05039_));
 sky130_fd_sc_hd__o22a_2 _24921_ (.A1(_05035_),
    .A2(_05036_),
    .B1(_05039_),
    .B2(_04997_),
    .X(_05040_));
 sky130_fd_sc_hd__clkbuf_2 _24922_ (.A(_05040_),
    .X(_05041_));
 sky130_fd_sc_hd__mux2_1 _24923_ (.A0(\cpuregs[4][5] ),
    .A1(_05041_),
    .S(_04994_),
    .X(_05042_));
 sky130_fd_sc_hd__clkbuf_1 _24924_ (.A(_05042_),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _24925_ (.A0(\reg_out[6] ),
    .A1(\alu_out_q[6] ),
    .S(_04979_),
    .X(_05043_));
 sky130_fd_sc_hd__and2_1 _24926_ (.A(_04978_),
    .B(_05043_),
    .X(_05044_));
 sky130_fd_sc_hd__clkbuf_2 _24927_ (.A(_04974_),
    .X(_05045_));
 sky130_fd_sc_hd__a221o_1 _24928_ (.A1(_05002_),
    .A2(\reg_next_pc[6] ),
    .B1(_08266_),
    .B2(_05003_),
    .C1(_05045_),
    .X(_05046_));
 sky130_fd_sc_hd__xor2_1 _24929_ (.A(_08997_),
    .B(_05037_),
    .X(_05047_));
 sky130_fd_sc_hd__o22a_4 _24930_ (.A1(_05044_),
    .A2(_05046_),
    .B1(_05047_),
    .B2(_04997_),
    .X(_05048_));
 sky130_fd_sc_hd__clkbuf_2 _24931_ (.A(_05048_),
    .X(_05049_));
 sky130_fd_sc_hd__clkbuf_4 _24932_ (.A(_04993_),
    .X(_05050_));
 sky130_fd_sc_hd__mux2_1 _24933_ (.A0(\cpuregs[4][6] ),
    .A1(_05049_),
    .S(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__clkbuf_1 _24934_ (.A(_05051_),
    .X(_00120_));
 sky130_fd_sc_hd__clkbuf_2 _24935_ (.A(_04972_),
    .X(_05052_));
 sky130_fd_sc_hd__mux2_1 _24936_ (.A0(\reg_out[7] ),
    .A1(\alu_out_q[7] ),
    .S(_04979_),
    .X(_05053_));
 sky130_fd_sc_hd__a221o_1 _24937_ (.A1(_05003_),
    .A2(_08273_),
    .B1(_04978_),
    .B2(_05053_),
    .C1(_05045_),
    .X(_05054_));
 sky130_fd_sc_hd__a21oi_1 _24938_ (.A1(_05052_),
    .A2(\reg_next_pc[7] ),
    .B1(_05054_),
    .Y(_05055_));
 sky130_fd_sc_hd__and3_1 _24939_ (.A(\reg_pc[7] ),
    .B(_08997_),
    .C(_05037_),
    .X(_05056_));
 sky130_fd_sc_hd__a21oi_1 _24940_ (.A1(_08997_),
    .A2(_05037_),
    .B1(\reg_pc[7] ),
    .Y(_05057_));
 sky130_fd_sc_hd__o21a_1 _24941_ (.A1(_05056_),
    .A2(_05057_),
    .B1(_05009_),
    .X(_05058_));
 sky130_fd_sc_hd__nor2_4 _24942_ (.A(_05055_),
    .B(_05058_),
    .Y(_05059_));
 sky130_fd_sc_hd__clkbuf_2 _24943_ (.A(_05059_),
    .X(_05060_));
 sky130_fd_sc_hd__mux2_1 _24944_ (.A0(\cpuregs[4][7] ),
    .A1(_05060_),
    .S(_05050_),
    .X(_05061_));
 sky130_fd_sc_hd__clkbuf_1 _24945_ (.A(_05061_),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _24946_ (.A0(\reg_out[8] ),
    .A1(\alu_out_q[8] ),
    .S(_04980_),
    .X(_05062_));
 sky130_fd_sc_hd__a221o_1 _24947_ (.A1(_05011_),
    .A2(_08237_),
    .B1(_04998_),
    .B2(_05062_),
    .C1(_05012_),
    .X(_05063_));
 sky130_fd_sc_hd__a21oi_1 _24948_ (.A1(_05052_),
    .A2(\reg_next_pc[8] ),
    .B1(_05063_),
    .Y(_05064_));
 sky130_fd_sc_hd__and2_1 _24949_ (.A(\reg_pc[8] ),
    .B(_05056_),
    .X(_05065_));
 sky130_fd_sc_hd__nor2_1 _24950_ (.A(\reg_pc[8] ),
    .B(_05056_),
    .Y(_05066_));
 sky130_fd_sc_hd__o21a_1 _24951_ (.A1(_05065_),
    .A2(_05066_),
    .B1(_05009_),
    .X(_05067_));
 sky130_fd_sc_hd__nor2_4 _24952_ (.A(_05064_),
    .B(_05067_),
    .Y(_05068_));
 sky130_fd_sc_hd__clkbuf_2 _24953_ (.A(_05068_),
    .X(_05069_));
 sky130_fd_sc_hd__mux2_1 _24954_ (.A0(\cpuregs[4][8] ),
    .A1(_05069_),
    .S(_05050_),
    .X(_05070_));
 sky130_fd_sc_hd__clkbuf_1 _24955_ (.A(_05070_),
    .X(_00122_));
 sky130_fd_sc_hd__xnor2_1 _24956_ (.A(_09170_),
    .B(_05065_),
    .Y(_05071_));
 sky130_fd_sc_hd__mux2_1 _24957_ (.A0(\reg_out[9] ),
    .A1(\alu_out_q[9] ),
    .S(_04980_),
    .X(_05072_));
 sky130_fd_sc_hd__a221o_1 _24958_ (.A1(_05011_),
    .A2(_08252_),
    .B1(_04998_),
    .B2(_05072_),
    .C1(_05012_),
    .X(_05073_));
 sky130_fd_sc_hd__a21oi_1 _24959_ (.A1(_04972_),
    .A2(\reg_next_pc[9] ),
    .B1(_05073_),
    .Y(_05074_));
 sky130_fd_sc_hd__a21oi_4 _24960_ (.A1(_05009_),
    .A2(_05071_),
    .B1(_05074_),
    .Y(_05075_));
 sky130_fd_sc_hd__clkbuf_2 _24961_ (.A(_05075_),
    .X(_05076_));
 sky130_fd_sc_hd__mux2_1 _24962_ (.A0(\cpuregs[4][9] ),
    .A1(_05076_),
    .S(_05050_),
    .X(_05077_));
 sky130_fd_sc_hd__clkbuf_1 _24963_ (.A(_05077_),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _24964_ (.A0(\reg_out[10] ),
    .A1(\alu_out_q[10] ),
    .S(_04980_),
    .X(_05078_));
 sky130_fd_sc_hd__a221o_1 _24965_ (.A1(_05011_),
    .A2(_08247_),
    .B1(_04998_),
    .B2(_05078_),
    .C1(_05012_),
    .X(_05079_));
 sky130_fd_sc_hd__a21oi_1 _24966_ (.A1(_05052_),
    .A2(\reg_next_pc[10] ),
    .B1(_05079_),
    .Y(_05080_));
 sky130_fd_sc_hd__and3_1 _24967_ (.A(_09218_),
    .B(_09170_),
    .C(_05065_),
    .X(_05081_));
 sky130_fd_sc_hd__a21oi_1 _24968_ (.A1(_09170_),
    .A2(_05065_),
    .B1(_09218_),
    .Y(_05082_));
 sky130_fd_sc_hd__o21a_1 _24969_ (.A1(_05081_),
    .A2(_05082_),
    .B1(_05009_),
    .X(_05083_));
 sky130_fd_sc_hd__nor2_4 _24970_ (.A(_05080_),
    .B(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__buf_2 _24971_ (.A(_05084_),
    .X(_05085_));
 sky130_fd_sc_hd__mux2_1 _24972_ (.A0(\cpuregs[4][10] ),
    .A1(_05085_),
    .S(_05050_),
    .X(_05086_));
 sky130_fd_sc_hd__clkbuf_1 _24973_ (.A(_05086_),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _24974_ (.A0(\reg_out[11] ),
    .A1(\alu_out_q[11] ),
    .S(_04980_),
    .X(_05087_));
 sky130_fd_sc_hd__a221o_1 _24975_ (.A1(_05011_),
    .A2(_08235_),
    .B1(_04998_),
    .B2(_05087_),
    .C1(_05012_),
    .X(_05088_));
 sky130_fd_sc_hd__a21oi_1 _24976_ (.A1(_05052_),
    .A2(\reg_next_pc[11] ),
    .B1(_05088_),
    .Y(_05089_));
 sky130_fd_sc_hd__and2_1 _24977_ (.A(_09295_),
    .B(_05081_),
    .X(_05090_));
 sky130_fd_sc_hd__nor2_1 _24978_ (.A(_09295_),
    .B(_05081_),
    .Y(_05091_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _24979_ (.A(_04974_),
    .X(_05092_));
 sky130_fd_sc_hd__o21a_1 _24980_ (.A1(_05090_),
    .A2(_05091_),
    .B1(_05092_),
    .X(_05093_));
 sky130_fd_sc_hd__nor2_4 _24981_ (.A(_05089_),
    .B(_05093_),
    .Y(_05094_));
 sky130_fd_sc_hd__clkbuf_2 _24982_ (.A(_05094_),
    .X(_05095_));
 sky130_fd_sc_hd__mux2_1 _24983_ (.A0(\cpuregs[4][11] ),
    .A1(_05095_),
    .S(_05050_),
    .X(_05096_));
 sky130_fd_sc_hd__clkbuf_1 _24984_ (.A(_05096_),
    .X(_00125_));
 sky130_fd_sc_hd__xnor2_1 _24985_ (.A(_09347_),
    .B(_05090_),
    .Y(_05097_));
 sky130_fd_sc_hd__mux2_1 _24986_ (.A0(\reg_out[12] ),
    .A1(\alu_out_q[12] ),
    .S(_04980_),
    .X(_05098_));
 sky130_fd_sc_hd__a221o_1 _24987_ (.A1(_05011_),
    .A2(_08251_),
    .B1(_04998_),
    .B2(_05098_),
    .C1(_05012_),
    .X(_05099_));
 sky130_fd_sc_hd__a21oi_1 _24988_ (.A1(_04972_),
    .A2(\reg_next_pc[12] ),
    .B1(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__a21oi_4 _24989_ (.A1(_05009_),
    .A2(_05097_),
    .B1(_05100_),
    .Y(_05101_));
 sky130_fd_sc_hd__clkbuf_2 _24990_ (.A(_05101_),
    .X(_05102_));
 sky130_fd_sc_hd__buf_2 _24991_ (.A(_04993_),
    .X(_05103_));
 sky130_fd_sc_hd__mux2_1 _24992_ (.A0(\cpuregs[4][12] ),
    .A1(_05102_),
    .S(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__clkbuf_1 _24993_ (.A(_05104_),
    .X(_00126_));
 sky130_fd_sc_hd__buf_2 _24994_ (.A(_04999_),
    .X(_05105_));
 sky130_fd_sc_hd__mux2_1 _24995_ (.A0(\reg_out[13] ),
    .A1(\alu_out_q[13] ),
    .S(_04981_),
    .X(_05106_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _24996_ (.A(_04971_),
    .X(_05107_));
 sky130_fd_sc_hd__a22o_1 _24997_ (.A1(_05107_),
    .A2(\reg_next_pc[13] ),
    .B1(_08260_),
    .B2(_10305_),
    .X(_05108_));
 sky130_fd_sc_hd__and3_1 _24998_ (.A(\reg_pc[13] ),
    .B(_09347_),
    .C(_05090_),
    .X(_05109_));
 sky130_fd_sc_hd__a31o_1 _24999_ (.A1(_09347_),
    .A2(_09295_),
    .A3(_05081_),
    .B1(\reg_pc[13] ),
    .X(_05110_));
 sky130_fd_sc_hd__and3b_1 _25000_ (.A_N(_05109_),
    .B(_05110_),
    .C(_05045_),
    .X(_05111_));
 sky130_fd_sc_hd__a211o_2 _25001_ (.A1(_05105_),
    .A2(_05106_),
    .B1(_05108_),
    .C1(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__clkbuf_2 _25002_ (.A(_05112_),
    .X(_05113_));
 sky130_fd_sc_hd__mux2_1 _25003_ (.A0(\cpuregs[4][13] ),
    .A1(_05113_),
    .S(_05103_),
    .X(_05114_));
 sky130_fd_sc_hd__clkbuf_1 _25004_ (.A(_05114_),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_1 _25005_ (.A0(\reg_out[14] ),
    .A1(\alu_out_q[14] ),
    .S(_04981_),
    .X(_05115_));
 sky130_fd_sc_hd__a22o_1 _25006_ (.A1(_05107_),
    .A2(\reg_next_pc[14] ),
    .B1(_08271_),
    .B2(_10305_),
    .X(_05116_));
 sky130_fd_sc_hd__and2_1 _25007_ (.A(_09386_),
    .B(_05109_),
    .X(_05117_));
 sky130_fd_sc_hd__o21ai_1 _25008_ (.A1(_09386_),
    .A2(_05109_),
    .B1(_05092_),
    .Y(_05118_));
 sky130_fd_sc_hd__nor2_1 _25009_ (.A(_05117_),
    .B(_05118_),
    .Y(_05119_));
 sky130_fd_sc_hd__a211o_2 _25010_ (.A1(_05105_),
    .A2(_05115_),
    .B1(_05116_),
    .C1(_05119_),
    .X(_05120_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _25011_ (.A(_05120_),
    .X(_05121_));
 sky130_fd_sc_hd__mux2_1 _25012_ (.A0(\cpuregs[4][14] ),
    .A1(_05121_),
    .S(_05103_),
    .X(_05122_));
 sky130_fd_sc_hd__clkbuf_1 _25013_ (.A(_05122_),
    .X(_00128_));
 sky130_fd_sc_hd__mux2_1 _25014_ (.A0(\reg_out[15] ),
    .A1(\alu_out_q[15] ),
    .S(_04981_),
    .X(_05123_));
 sky130_fd_sc_hd__a22o_1 _25015_ (.A1(_05107_),
    .A2(\reg_next_pc[15] ),
    .B1(_08250_),
    .B2(_10305_),
    .X(_05124_));
 sky130_fd_sc_hd__and3_1 _25016_ (.A(\reg_pc[15] ),
    .B(_09386_),
    .C(_05109_),
    .X(_05125_));
 sky130_fd_sc_hd__o21ai_1 _25017_ (.A1(\reg_pc[15] ),
    .A2(_05117_),
    .B1(_05092_),
    .Y(_05126_));
 sky130_fd_sc_hd__nor2_1 _25018_ (.A(_05125_),
    .B(_05126_),
    .Y(_05127_));
 sky130_fd_sc_hd__a211o_4 _25019_ (.A1(_05105_),
    .A2(_05123_),
    .B1(_05124_),
    .C1(_05127_),
    .X(_05128_));
 sky130_fd_sc_hd__clkbuf_2 _25020_ (.A(_05128_),
    .X(_05129_));
 sky130_fd_sc_hd__mux2_1 _25021_ (.A0(\cpuregs[4][15] ),
    .A1(_05129_),
    .S(_05103_),
    .X(_05130_));
 sky130_fd_sc_hd__clkbuf_1 _25022_ (.A(_05130_),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_1 _25023_ (.A0(\reg_out[16] ),
    .A1(\alu_out_q[16] ),
    .S(_04981_),
    .X(_05131_));
 sky130_fd_sc_hd__clkbuf_2 _25024_ (.A(_10304_),
    .X(_05132_));
 sky130_fd_sc_hd__a22o_1 _25025_ (.A1(_05107_),
    .A2(\reg_next_pc[16] ),
    .B1(_08257_),
    .B2(_05132_),
    .X(_05133_));
 sky130_fd_sc_hd__and2_1 _25026_ (.A(_09468_),
    .B(_05125_),
    .X(_05134_));
 sky130_fd_sc_hd__o21ai_1 _25027_ (.A1(_09468_),
    .A2(_05125_),
    .B1(_05092_),
    .Y(_05135_));
 sky130_fd_sc_hd__nor2_1 _25028_ (.A(_05134_),
    .B(_05135_),
    .Y(_05136_));
 sky130_fd_sc_hd__a211o_4 _25029_ (.A1(_05105_),
    .A2(_05131_),
    .B1(_05133_),
    .C1(_05136_),
    .X(_05137_));
 sky130_fd_sc_hd__clkbuf_2 _25030_ (.A(_05137_),
    .X(_05138_));
 sky130_fd_sc_hd__mux2_1 _25031_ (.A0(\cpuregs[4][16] ),
    .A1(_05138_),
    .S(_05103_),
    .X(_05139_));
 sky130_fd_sc_hd__clkbuf_1 _25032_ (.A(_05139_),
    .X(_00130_));
 sky130_fd_sc_hd__mux2_1 _25033_ (.A0(\reg_out[17] ),
    .A1(\alu_out_q[17] ),
    .S(_04981_),
    .X(_05140_));
 sky130_fd_sc_hd__a22o_1 _25034_ (.A1(_05107_),
    .A2(\reg_next_pc[17] ),
    .B1(_08272_),
    .B2(_05132_),
    .X(_05141_));
 sky130_fd_sc_hd__and3_1 _25035_ (.A(\reg_pc[17] ),
    .B(_09468_),
    .C(_05125_),
    .X(_05142_));
 sky130_fd_sc_hd__o21ai_1 _25036_ (.A1(\reg_pc[17] ),
    .A2(_05134_),
    .B1(_05092_),
    .Y(_05143_));
 sky130_fd_sc_hd__nor2_1 _25037_ (.A(_05142_),
    .B(_05143_),
    .Y(_05144_));
 sky130_fd_sc_hd__a211o_4 _25038_ (.A1(_05105_),
    .A2(_05140_),
    .B1(_05141_),
    .C1(_05144_),
    .X(_05145_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _25039_ (.A(_05145_),
    .X(_05146_));
 sky130_fd_sc_hd__mux2_1 _25040_ (.A0(\cpuregs[4][17] ),
    .A1(_05146_),
    .S(_05103_),
    .X(_05147_));
 sky130_fd_sc_hd__clkbuf_1 _25041_ (.A(_05147_),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_2 _25042_ (.A0(\reg_out[18] ),
    .A1(\alu_out_q[18] ),
    .S(_04982_),
    .X(_05148_));
 sky130_fd_sc_hd__a22o_1 _25043_ (.A1(_05107_),
    .A2(\reg_next_pc[18] ),
    .B1(_08234_),
    .B2(_05132_),
    .X(_05149_));
 sky130_fd_sc_hd__clkbuf_2 _25044_ (.A(\reg_pc[18] ),
    .X(_05150_));
 sky130_fd_sc_hd__a21oi_1 _25045_ (.A1(_05150_),
    .A2(_05142_),
    .B1(_04997_),
    .Y(_05151_));
 sky130_fd_sc_hd__o21a_1 _25046_ (.A1(_05150_),
    .A2(_05142_),
    .B1(_05151_),
    .X(_05152_));
 sky130_fd_sc_hd__a211o_4 _25047_ (.A1(_05105_),
    .A2(_05148_),
    .B1(_05149_),
    .C1(_05152_),
    .X(_05153_));
 sky130_fd_sc_hd__clkbuf_2 _25048_ (.A(_05153_),
    .X(_05154_));
 sky130_fd_sc_hd__buf_2 _25049_ (.A(_04993_),
    .X(_05155_));
 sky130_fd_sc_hd__mux2_1 _25050_ (.A0(\cpuregs[4][18] ),
    .A1(_05154_),
    .S(_05155_),
    .X(_05156_));
 sky130_fd_sc_hd__clkbuf_1 _25051_ (.A(_05156_),
    .X(_00132_));
 sky130_fd_sc_hd__buf_2 _25052_ (.A(_04999_),
    .X(_05157_));
 sky130_fd_sc_hd__mux2_2 _25053_ (.A0(\reg_out[19] ),
    .A1(\alu_out_q[19] ),
    .S(_04982_),
    .X(_05158_));
 sky130_fd_sc_hd__clkbuf_2 _25054_ (.A(_04971_),
    .X(_05159_));
 sky130_fd_sc_hd__a22o_1 _25055_ (.A1(_05159_),
    .A2(\reg_next_pc[19] ),
    .B1(_08255_),
    .B2(_05132_),
    .X(_05160_));
 sky130_fd_sc_hd__and3_1 _25056_ (.A(\reg_pc[19] ),
    .B(_05150_),
    .C(_05142_),
    .X(_05161_));
 sky130_fd_sc_hd__a21o_1 _25057_ (.A1(_05150_),
    .A2(_05142_),
    .B1(\reg_pc[19] ),
    .X(_05162_));
 sky130_fd_sc_hd__and3b_1 _25058_ (.A_N(_05161_),
    .B(_05045_),
    .C(_05162_),
    .X(_05163_));
 sky130_fd_sc_hd__a211o_4 _25059_ (.A1(_05157_),
    .A2(_05158_),
    .B1(_05160_),
    .C1(_05163_),
    .X(_05164_));
 sky130_fd_sc_hd__buf_2 _25060_ (.A(_05164_),
    .X(_05165_));
 sky130_fd_sc_hd__mux2_1 _25061_ (.A0(\cpuregs[4][19] ),
    .A1(_05165_),
    .S(_05155_),
    .X(_05166_));
 sky130_fd_sc_hd__clkbuf_1 _25062_ (.A(_05166_),
    .X(_00133_));
 sky130_fd_sc_hd__mux2_2 _25063_ (.A0(\reg_out[20] ),
    .A1(\alu_out_q[20] ),
    .S(_04982_),
    .X(_05167_));
 sky130_fd_sc_hd__a22o_1 _25064_ (.A1(_05159_),
    .A2(\reg_next_pc[20] ),
    .B1(_08244_),
    .B2(_05132_),
    .X(_05168_));
 sky130_fd_sc_hd__and2_1 _25065_ (.A(_09634_),
    .B(_05161_),
    .X(_05169_));
 sky130_fd_sc_hd__o21ai_1 _25066_ (.A1(_09634_),
    .A2(_05161_),
    .B1(_05092_),
    .Y(_05170_));
 sky130_fd_sc_hd__nor2_1 _25067_ (.A(_05169_),
    .B(_05170_),
    .Y(_05171_));
 sky130_fd_sc_hd__a211o_4 _25068_ (.A1(_05157_),
    .A2(_05167_),
    .B1(_05168_),
    .C1(_05171_),
    .X(_05172_));
 sky130_fd_sc_hd__clkbuf_2 _25069_ (.A(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__mux2_1 _25070_ (.A0(\cpuregs[4][20] ),
    .A1(_05173_),
    .S(_05155_),
    .X(_05174_));
 sky130_fd_sc_hd__clkbuf_1 _25071_ (.A(_05174_),
    .X(_00134_));
 sky130_fd_sc_hd__mux2_2 _25072_ (.A0(\reg_out[21] ),
    .A1(\alu_out_q[21] ),
    .S(_04982_),
    .X(_05175_));
 sky130_fd_sc_hd__a22o_1 _25073_ (.A1(_05159_),
    .A2(\reg_next_pc[21] ),
    .B1(_08246_),
    .B2(_05132_),
    .X(_05176_));
 sky130_fd_sc_hd__and3_1 _25074_ (.A(\reg_pc[21] ),
    .B(_09634_),
    .C(_05161_),
    .X(_05177_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _25075_ (.A(_04974_),
    .X(_05178_));
 sky130_fd_sc_hd__o21ai_1 _25076_ (.A1(\reg_pc[21] ),
    .A2(_05169_),
    .B1(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hd__nor2_1 _25077_ (.A(_05177_),
    .B(_05179_),
    .Y(_05180_));
 sky130_fd_sc_hd__a211o_4 _25078_ (.A1(_05157_),
    .A2(_05175_),
    .B1(_05176_),
    .C1(_05180_),
    .X(_05181_));
 sky130_fd_sc_hd__buf_2 _25079_ (.A(_05181_),
    .X(_05182_));
 sky130_fd_sc_hd__mux2_1 _25080_ (.A0(\cpuregs[4][21] ),
    .A1(_05182_),
    .S(_05155_),
    .X(_05183_));
 sky130_fd_sc_hd__clkbuf_1 _25081_ (.A(_05183_),
    .X(_00135_));
 sky130_fd_sc_hd__mux2_2 _25082_ (.A0(\reg_out[22] ),
    .A1(\alu_out_q[22] ),
    .S(_04982_),
    .X(_05184_));
 sky130_fd_sc_hd__clkbuf_2 _25083_ (.A(_10304_),
    .X(_05185_));
 sky130_fd_sc_hd__a22o_1 _25084_ (.A1(_05159_),
    .A2(\reg_next_pc[22] ),
    .B1(_08245_),
    .B2(_05185_),
    .X(_05186_));
 sky130_fd_sc_hd__and2_1 _25085_ (.A(_09712_),
    .B(_05177_),
    .X(_05187_));
 sky130_fd_sc_hd__o21ai_1 _25086_ (.A1(_09712_),
    .A2(_05177_),
    .B1(_05178_),
    .Y(_05188_));
 sky130_fd_sc_hd__nor2_1 _25087_ (.A(_05187_),
    .B(_05188_),
    .Y(_05189_));
 sky130_fd_sc_hd__a211o_4 _25088_ (.A1(_05157_),
    .A2(_05184_),
    .B1(_05186_),
    .C1(_05189_),
    .X(_05190_));
 sky130_fd_sc_hd__buf_2 _25089_ (.A(_05190_),
    .X(_05191_));
 sky130_fd_sc_hd__mux2_1 _25090_ (.A0(\cpuregs[4][22] ),
    .A1(_05191_),
    .S(_05155_),
    .X(_05192_));
 sky130_fd_sc_hd__clkbuf_1 _25091_ (.A(_05192_),
    .X(_00136_));
 sky130_fd_sc_hd__mux2_1 _25092_ (.A0(\reg_out[23] ),
    .A1(\alu_out_q[23] ),
    .S(_04983_),
    .X(_05193_));
 sky130_fd_sc_hd__a22o_1 _25093_ (.A1(_05159_),
    .A2(\reg_next_pc[23] ),
    .B1(_08249_),
    .B2(_05185_),
    .X(_05194_));
 sky130_fd_sc_hd__and3_1 _25094_ (.A(\reg_pc[23] ),
    .B(_09712_),
    .C(_05177_),
    .X(_05195_));
 sky130_fd_sc_hd__o21ai_1 _25095_ (.A1(_09750_),
    .A2(_05187_),
    .B1(_05178_),
    .Y(_05196_));
 sky130_fd_sc_hd__nor2_1 _25096_ (.A(_05195_),
    .B(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__a211o_4 _25097_ (.A1(_05157_),
    .A2(_05193_),
    .B1(_05194_),
    .C1(_05197_),
    .X(_05198_));
 sky130_fd_sc_hd__clkbuf_2 _25098_ (.A(_05198_),
    .X(_05199_));
 sky130_fd_sc_hd__mux2_1 _25099_ (.A0(\cpuregs[4][23] ),
    .A1(_05199_),
    .S(_05155_),
    .X(_05200_));
 sky130_fd_sc_hd__clkbuf_1 _25100_ (.A(_05200_),
    .X(_00137_));
 sky130_fd_sc_hd__mux2_1 _25101_ (.A0(\reg_out[24] ),
    .A1(\alu_out_q[24] ),
    .S(_04983_),
    .X(_05201_));
 sky130_fd_sc_hd__a22o_1 _25102_ (.A1(_05159_),
    .A2(\reg_next_pc[24] ),
    .B1(_08262_),
    .B2(_05185_),
    .X(_05202_));
 sky130_fd_sc_hd__a21oi_1 _25103_ (.A1(_09788_),
    .A2(_05195_),
    .B1(_04996_),
    .Y(_05203_));
 sky130_fd_sc_hd__o21a_1 _25104_ (.A1(_09788_),
    .A2(_05195_),
    .B1(_05203_),
    .X(_05204_));
 sky130_fd_sc_hd__a211o_4 _25105_ (.A1(_05157_),
    .A2(_05201_),
    .B1(_05202_),
    .C1(_05204_),
    .X(_05205_));
 sky130_fd_sc_hd__clkbuf_2 _25106_ (.A(_05205_),
    .X(_05206_));
 sky130_fd_sc_hd__buf_2 _25107_ (.A(_04992_),
    .X(_05207_));
 sky130_fd_sc_hd__mux2_1 _25108_ (.A0(\cpuregs[4][24] ),
    .A1(_05206_),
    .S(_05207_),
    .X(_05208_));
 sky130_fd_sc_hd__clkbuf_1 _25109_ (.A(_05208_),
    .X(_00138_));
 sky130_fd_sc_hd__buf_2 _25110_ (.A(_04999_),
    .X(_05209_));
 sky130_fd_sc_hd__mux2_1 _25111_ (.A0(\reg_out[25] ),
    .A1(\alu_out_q[25] ),
    .S(_04983_),
    .X(_05210_));
 sky130_fd_sc_hd__clkbuf_2 _25112_ (.A(_04971_),
    .X(_05211_));
 sky130_fd_sc_hd__a22o_1 _25113_ (.A1(_05211_),
    .A2(\reg_next_pc[25] ),
    .B1(_08239_),
    .B2(_05185_),
    .X(_05212_));
 sky130_fd_sc_hd__and3_1 _25114_ (.A(\reg_pc[25] ),
    .B(\reg_pc[24] ),
    .C(_05195_),
    .X(_05213_));
 sky130_fd_sc_hd__a21o_1 _25115_ (.A1(_09788_),
    .A2(_05195_),
    .B1(\reg_pc[25] ),
    .X(_05214_));
 sky130_fd_sc_hd__and3b_1 _25116_ (.A_N(_05213_),
    .B(_05045_),
    .C(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__a211o_4 _25117_ (.A1(_05209_),
    .A2(_05210_),
    .B1(_05212_),
    .C1(_05215_),
    .X(_05216_));
 sky130_fd_sc_hd__clkbuf_2 _25118_ (.A(_05216_),
    .X(_05217_));
 sky130_fd_sc_hd__mux2_1 _25119_ (.A0(\cpuregs[4][25] ),
    .A1(_05217_),
    .S(_05207_),
    .X(_05218_));
 sky130_fd_sc_hd__clkbuf_1 _25120_ (.A(_05218_),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_1 _25121_ (.A0(\reg_out[26] ),
    .A1(\alu_out_q[26] ),
    .S(_04983_),
    .X(_05219_));
 sky130_fd_sc_hd__a22o_1 _25122_ (.A1(_05211_),
    .A2(\reg_next_pc[26] ),
    .B1(_08241_),
    .B2(_05185_),
    .X(_05220_));
 sky130_fd_sc_hd__and2_1 _25123_ (.A(\reg_pc[26] ),
    .B(_05213_),
    .X(_05221_));
 sky130_fd_sc_hd__o21ai_1 _25124_ (.A1(_09894_),
    .A2(_05213_),
    .B1(_05178_),
    .Y(_05222_));
 sky130_fd_sc_hd__nor2_1 _25125_ (.A(_05221_),
    .B(_05222_),
    .Y(_05223_));
 sky130_fd_sc_hd__a211o_4 _25126_ (.A1(_05209_),
    .A2(_05219_),
    .B1(_05220_),
    .C1(_05223_),
    .X(_05224_));
 sky130_fd_sc_hd__clkbuf_2 _25127_ (.A(_05224_),
    .X(_05225_));
 sky130_fd_sc_hd__mux2_1 _25128_ (.A0(\cpuregs[4][26] ),
    .A1(_05225_),
    .S(_05207_),
    .X(_05226_));
 sky130_fd_sc_hd__clkbuf_1 _25129_ (.A(_05226_),
    .X(_00140_));
 sky130_fd_sc_hd__mux2_1 _25130_ (.A0(\reg_out[27] ),
    .A1(\alu_out_q[27] ),
    .S(_04984_),
    .X(_05227_));
 sky130_fd_sc_hd__a22o_1 _25131_ (.A1(_05211_),
    .A2(\reg_next_pc[27] ),
    .B1(_08261_),
    .B2(_05185_),
    .X(_05228_));
 sky130_fd_sc_hd__a21oi_1 _25132_ (.A1(_09902_),
    .A2(_05221_),
    .B1(_04996_),
    .Y(_05229_));
 sky130_fd_sc_hd__o21a_1 _25133_ (.A1(_09902_),
    .A2(_05221_),
    .B1(_05229_),
    .X(_05230_));
 sky130_fd_sc_hd__a211o_4 _25134_ (.A1(_05209_),
    .A2(_05227_),
    .B1(_05228_),
    .C1(_05230_),
    .X(_05231_));
 sky130_fd_sc_hd__clkbuf_2 _25135_ (.A(_05231_),
    .X(_05232_));
 sky130_fd_sc_hd__mux2_1 _25136_ (.A0(\cpuregs[4][27] ),
    .A1(_05232_),
    .S(_05207_),
    .X(_05233_));
 sky130_fd_sc_hd__clkbuf_1 _25137_ (.A(_05233_),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_1 _25138_ (.A0(\reg_out[28] ),
    .A1(\alu_out_q[28] ),
    .S(_04983_),
    .X(_05234_));
 sky130_fd_sc_hd__a22o_1 _25139_ (.A1(_05211_),
    .A2(\reg_next_pc[28] ),
    .B1(_08256_),
    .B2(_04977_),
    .X(_05235_));
 sky130_fd_sc_hd__and3_1 _25140_ (.A(\reg_pc[28] ),
    .B(\reg_pc[27] ),
    .C(_05221_),
    .X(_05236_));
 sky130_fd_sc_hd__a31o_1 _25141_ (.A1(_09902_),
    .A2(_09894_),
    .A3(_05213_),
    .B1(\reg_pc[28] ),
    .X(_05237_));
 sky130_fd_sc_hd__and3b_1 _25142_ (.A_N(_05236_),
    .B(_05237_),
    .C(_05045_),
    .X(_05238_));
 sky130_fd_sc_hd__a211o_4 _25143_ (.A1(_05209_),
    .A2(_05234_),
    .B1(_05235_),
    .C1(_05238_),
    .X(_05239_));
 sky130_fd_sc_hd__clkbuf_2 _25144_ (.A(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__mux2_1 _25145_ (.A0(\cpuregs[4][28] ),
    .A1(_05240_),
    .S(_05207_),
    .X(_05241_));
 sky130_fd_sc_hd__clkbuf_1 _25146_ (.A(_05241_),
    .X(_00142_));
 sky130_fd_sc_hd__mux2_1 _25147_ (.A0(\reg_out[29] ),
    .A1(\alu_out_q[29] ),
    .S(_04984_),
    .X(_05242_));
 sky130_fd_sc_hd__a22o_1 _25148_ (.A1(_05211_),
    .A2(\reg_next_pc[29] ),
    .B1(_08242_),
    .B2(_04977_),
    .X(_05243_));
 sky130_fd_sc_hd__and2_1 _25149_ (.A(_09975_),
    .B(_05236_),
    .X(_05244_));
 sky130_fd_sc_hd__o21ai_1 _25150_ (.A1(_09975_),
    .A2(_05236_),
    .B1(_05178_),
    .Y(_05245_));
 sky130_fd_sc_hd__nor2_1 _25151_ (.A(_05244_),
    .B(_05245_),
    .Y(_05246_));
 sky130_fd_sc_hd__a211o_4 _25152_ (.A1(_05209_),
    .A2(_05242_),
    .B1(_05243_),
    .C1(_05246_),
    .X(_05247_));
 sky130_fd_sc_hd__clkbuf_2 _25153_ (.A(_05247_),
    .X(_05248_));
 sky130_fd_sc_hd__mux2_1 _25154_ (.A0(\cpuregs[4][29] ),
    .A1(_05248_),
    .S(_05207_),
    .X(_05249_));
 sky130_fd_sc_hd__clkbuf_1 _25155_ (.A(_05249_),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _25156_ (.A0(\reg_out[30] ),
    .A1(\alu_out_q[30] ),
    .S(_04984_),
    .X(_05250_));
 sky130_fd_sc_hd__a22o_1 _25157_ (.A1(_05211_),
    .A2(\reg_next_pc[30] ),
    .B1(_08270_),
    .B2(_04977_),
    .X(_05251_));
 sky130_fd_sc_hd__and3_1 _25158_ (.A(\reg_pc[30] ),
    .B(\reg_pc[29] ),
    .C(_05236_),
    .X(_05252_));
 sky130_fd_sc_hd__o21ai_1 _25159_ (.A1(\reg_pc[30] ),
    .A2(_05244_),
    .B1(_05178_),
    .Y(_05253_));
 sky130_fd_sc_hd__nor2_1 _25160_ (.A(_05252_),
    .B(_05253_),
    .Y(_05254_));
 sky130_fd_sc_hd__a211o_4 _25161_ (.A1(_05209_),
    .A2(_05250_),
    .B1(_05251_),
    .C1(_05254_),
    .X(_05255_));
 sky130_fd_sc_hd__clkbuf_2 _25162_ (.A(_05255_),
    .X(_05256_));
 sky130_fd_sc_hd__mux2_1 _25163_ (.A0(\cpuregs[4][30] ),
    .A1(_05256_),
    .S(_04993_),
    .X(_05257_));
 sky130_fd_sc_hd__clkbuf_1 _25164_ (.A(_05257_),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _25165_ (.A0(\reg_out[31] ),
    .A1(\alu_out_q[31] ),
    .S(_04984_),
    .X(_05258_));
 sky130_fd_sc_hd__a22o_1 _25166_ (.A1(_05002_),
    .A2(\reg_next_pc[31] ),
    .B1(_08258_),
    .B2(_04977_),
    .X(_05259_));
 sky130_fd_sc_hd__o21ai_1 _25167_ (.A1(\reg_pc[31] ),
    .A2(_05252_),
    .B1(_04975_),
    .Y(_05260_));
 sky130_fd_sc_hd__a21oi_1 _25168_ (.A1(\reg_pc[31] ),
    .A2(_05252_),
    .B1(_05260_),
    .Y(_05261_));
 sky130_fd_sc_hd__a211o_4 _25169_ (.A1(_04999_),
    .A2(_05258_),
    .B1(_05259_),
    .C1(_05261_),
    .X(_05262_));
 sky130_fd_sc_hd__buf_2 _25170_ (.A(_05262_),
    .X(_05263_));
 sky130_fd_sc_hd__mux2_1 _25171_ (.A0(\cpuregs[4][31] ),
    .A1(_05263_),
    .S(_04993_),
    .X(_05264_));
 sky130_fd_sc_hd__clkbuf_1 _25172_ (.A(_05264_),
    .X(_00145_));
 sky130_fd_sc_hd__buf_1 _25173_ (.A(_04987_),
    .X(_05265_));
 sky130_vsdinv _25174_ (.A(\latched_rd[1] ),
    .Y(_05266_));
 sky130_vsdinv _25175_ (.A(\latched_rd[0] ),
    .Y(_05267_));
 sky130_fd_sc_hd__or3_2 _25176_ (.A(_05266_),
    .B(_05267_),
    .C(_04989_),
    .X(_05268_));
 sky130_fd_sc_hd__or3_1 _25177_ (.A(\latched_rd[2] ),
    .B(\latched_rd[4] ),
    .C(\latched_rd[3] ),
    .X(_05269_));
 sky130_fd_sc_hd__or2_1 _25178_ (.A(_05268_),
    .B(_05269_),
    .X(_05270_));
 sky130_fd_sc_hd__buf_4 _25179_ (.A(_05270_),
    .X(_05271_));
 sky130_fd_sc_hd__buf_2 _25180_ (.A(_05271_),
    .X(_05272_));
 sky130_fd_sc_hd__mux2_1 _25181_ (.A0(_05265_),
    .A1(\cpuregs[3][0] ),
    .S(_05272_),
    .X(_05273_));
 sky130_fd_sc_hd__clkbuf_1 _25182_ (.A(_05273_),
    .X(_00146_));
 sky130_fd_sc_hd__clkbuf_2 _25183_ (.A(_05005_),
    .X(_05274_));
 sky130_fd_sc_hd__mux2_1 _25184_ (.A0(_05274_),
    .A1(\cpuregs[3][1] ),
    .S(_05272_),
    .X(_05275_));
 sky130_fd_sc_hd__clkbuf_1 _25185_ (.A(_05275_),
    .X(_00147_));
 sky130_fd_sc_hd__clkbuf_2 _25186_ (.A(_05015_),
    .X(_05276_));
 sky130_fd_sc_hd__mux2_1 _25187_ (.A0(_05276_),
    .A1(\cpuregs[3][2] ),
    .S(_05272_),
    .X(_05277_));
 sky130_fd_sc_hd__clkbuf_1 _25188_ (.A(_05277_),
    .X(_00148_));
 sky130_fd_sc_hd__clkbuf_2 _25189_ (.A(_05022_),
    .X(_05278_));
 sky130_fd_sc_hd__mux2_1 _25190_ (.A0(_05278_),
    .A1(\cpuregs[3][3] ),
    .S(_05272_),
    .X(_05279_));
 sky130_fd_sc_hd__clkbuf_1 _25191_ (.A(_05279_),
    .X(_00149_));
 sky130_fd_sc_hd__buf_1 _25192_ (.A(_05031_),
    .X(_05280_));
 sky130_fd_sc_hd__mux2_1 _25193_ (.A0(_05280_),
    .A1(\cpuregs[3][4] ),
    .S(_05272_),
    .X(_05281_));
 sky130_fd_sc_hd__clkbuf_1 _25194_ (.A(_05281_),
    .X(_00150_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _25195_ (.A(_05040_),
    .X(_05282_));
 sky130_fd_sc_hd__mux2_1 _25196_ (.A0(_05282_),
    .A1(\cpuregs[3][5] ),
    .S(_05272_),
    .X(_05283_));
 sky130_fd_sc_hd__clkbuf_1 _25197_ (.A(_05283_),
    .X(_00151_));
 sky130_fd_sc_hd__buf_1 _25198_ (.A(_05048_),
    .X(_05284_));
 sky130_fd_sc_hd__clkbuf_4 _25199_ (.A(_05271_),
    .X(_05285_));
 sky130_fd_sc_hd__mux2_1 _25200_ (.A0(_05284_),
    .A1(\cpuregs[3][6] ),
    .S(_05285_),
    .X(_05286_));
 sky130_fd_sc_hd__clkbuf_1 _25201_ (.A(_05286_),
    .X(_00152_));
 sky130_fd_sc_hd__buf_1 _25202_ (.A(_05059_),
    .X(_05287_));
 sky130_fd_sc_hd__mux2_1 _25203_ (.A0(_05287_),
    .A1(\cpuregs[3][7] ),
    .S(_05285_),
    .X(_05288_));
 sky130_fd_sc_hd__clkbuf_1 _25204_ (.A(_05288_),
    .X(_00153_));
 sky130_fd_sc_hd__buf_1 _25205_ (.A(_05068_),
    .X(_05289_));
 sky130_fd_sc_hd__mux2_1 _25206_ (.A0(_05289_),
    .A1(\cpuregs[3][8] ),
    .S(_05285_),
    .X(_05290_));
 sky130_fd_sc_hd__clkbuf_1 _25207_ (.A(_05290_),
    .X(_00154_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _25208_ (.A(_05075_),
    .X(_05291_));
 sky130_fd_sc_hd__mux2_1 _25209_ (.A0(_05291_),
    .A1(\cpuregs[3][9] ),
    .S(_05285_),
    .X(_05292_));
 sky130_fd_sc_hd__clkbuf_1 _25210_ (.A(_05292_),
    .X(_00155_));
 sky130_fd_sc_hd__buf_1 _25211_ (.A(_05084_),
    .X(_05293_));
 sky130_fd_sc_hd__mux2_1 _25212_ (.A0(_05293_),
    .A1(\cpuregs[3][10] ),
    .S(_05285_),
    .X(_05294_));
 sky130_fd_sc_hd__clkbuf_1 _25213_ (.A(_05294_),
    .X(_00156_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _25214_ (.A(_05094_),
    .X(_05295_));
 sky130_fd_sc_hd__mux2_1 _25215_ (.A0(_05295_),
    .A1(\cpuregs[3][11] ),
    .S(_05285_),
    .X(_05296_));
 sky130_fd_sc_hd__clkbuf_1 _25216_ (.A(_05296_),
    .X(_00157_));
 sky130_fd_sc_hd__clkbuf_2 _25217_ (.A(_05101_),
    .X(_05297_));
 sky130_fd_sc_hd__clkbuf_4 _25218_ (.A(_05271_),
    .X(_05298_));
 sky130_fd_sc_hd__mux2_1 _25219_ (.A0(_05297_),
    .A1(\cpuregs[3][12] ),
    .S(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__clkbuf_1 _25220_ (.A(_05299_),
    .X(_00158_));
 sky130_fd_sc_hd__clkbuf_2 _25221_ (.A(_05112_),
    .X(_05300_));
 sky130_fd_sc_hd__mux2_1 _25222_ (.A0(_05300_),
    .A1(\cpuregs[3][13] ),
    .S(_05298_),
    .X(_05301_));
 sky130_fd_sc_hd__clkbuf_1 _25223_ (.A(_05301_),
    .X(_00159_));
 sky130_fd_sc_hd__buf_2 _25224_ (.A(_05120_),
    .X(_05302_));
 sky130_fd_sc_hd__mux2_1 _25225_ (.A0(_05302_),
    .A1(\cpuregs[3][14] ),
    .S(_05298_),
    .X(_05303_));
 sky130_fd_sc_hd__clkbuf_1 _25226_ (.A(_05303_),
    .X(_00160_));
 sky130_fd_sc_hd__clkbuf_2 _25227_ (.A(_05128_),
    .X(_05304_));
 sky130_fd_sc_hd__mux2_1 _25228_ (.A0(_05304_),
    .A1(\cpuregs[3][15] ),
    .S(_05298_),
    .X(_05305_));
 sky130_fd_sc_hd__clkbuf_1 _25229_ (.A(_05305_),
    .X(_00161_));
 sky130_fd_sc_hd__clkbuf_2 _25230_ (.A(_05137_),
    .X(_05306_));
 sky130_fd_sc_hd__mux2_1 _25231_ (.A0(_05306_),
    .A1(\cpuregs[3][16] ),
    .S(_05298_),
    .X(_05307_));
 sky130_fd_sc_hd__clkbuf_1 _25232_ (.A(_05307_),
    .X(_00162_));
 sky130_fd_sc_hd__clkbuf_2 _25233_ (.A(_05145_),
    .X(_05308_));
 sky130_fd_sc_hd__mux2_1 _25234_ (.A0(_05308_),
    .A1(\cpuregs[3][17] ),
    .S(_05298_),
    .X(_05309_));
 sky130_fd_sc_hd__clkbuf_1 _25235_ (.A(_05309_),
    .X(_00163_));
 sky130_fd_sc_hd__clkbuf_2 _25236_ (.A(_05153_),
    .X(_05310_));
 sky130_fd_sc_hd__clkbuf_2 _25237_ (.A(_05271_),
    .X(_05311_));
 sky130_fd_sc_hd__mux2_1 _25238_ (.A0(_05310_),
    .A1(\cpuregs[3][18] ),
    .S(_05311_),
    .X(_05312_));
 sky130_fd_sc_hd__clkbuf_1 _25239_ (.A(_05312_),
    .X(_00164_));
 sky130_fd_sc_hd__clkbuf_2 _25240_ (.A(_05164_),
    .X(_05313_));
 sky130_fd_sc_hd__mux2_1 _25241_ (.A0(_05313_),
    .A1(\cpuregs[3][19] ),
    .S(_05311_),
    .X(_05314_));
 sky130_fd_sc_hd__clkbuf_1 _25242_ (.A(_05314_),
    .X(_00165_));
 sky130_fd_sc_hd__clkbuf_2 _25243_ (.A(_05172_),
    .X(_05315_));
 sky130_fd_sc_hd__mux2_1 _25244_ (.A0(_05315_),
    .A1(\cpuregs[3][20] ),
    .S(_05311_),
    .X(_05316_));
 sky130_fd_sc_hd__clkbuf_1 _25245_ (.A(_05316_),
    .X(_00166_));
 sky130_fd_sc_hd__clkbuf_2 _25246_ (.A(_05181_),
    .X(_05317_));
 sky130_fd_sc_hd__mux2_1 _25247_ (.A0(_05317_),
    .A1(\cpuregs[3][21] ),
    .S(_05311_),
    .X(_05318_));
 sky130_fd_sc_hd__clkbuf_1 _25248_ (.A(_05318_),
    .X(_00167_));
 sky130_fd_sc_hd__clkbuf_2 _25249_ (.A(_05190_),
    .X(_05319_));
 sky130_fd_sc_hd__mux2_1 _25250_ (.A0(_05319_),
    .A1(\cpuregs[3][22] ),
    .S(_05311_),
    .X(_05320_));
 sky130_fd_sc_hd__clkbuf_1 _25251_ (.A(_05320_),
    .X(_00168_));
 sky130_fd_sc_hd__clkbuf_2 _25252_ (.A(_05198_),
    .X(_05321_));
 sky130_fd_sc_hd__mux2_1 _25253_ (.A0(_05321_),
    .A1(\cpuregs[3][23] ),
    .S(_05311_),
    .X(_05322_));
 sky130_fd_sc_hd__clkbuf_1 _25254_ (.A(_05322_),
    .X(_00169_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _25255_ (.A(_05205_),
    .X(_05323_));
 sky130_fd_sc_hd__clkbuf_4 _25256_ (.A(_05270_),
    .X(_05324_));
 sky130_fd_sc_hd__mux2_1 _25257_ (.A0(_05323_),
    .A1(\cpuregs[3][24] ),
    .S(_05324_),
    .X(_05325_));
 sky130_fd_sc_hd__clkbuf_1 _25258_ (.A(_05325_),
    .X(_00170_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _25259_ (.A(_05216_),
    .X(_05326_));
 sky130_fd_sc_hd__mux2_1 _25260_ (.A0(_05326_),
    .A1(\cpuregs[3][25] ),
    .S(_05324_),
    .X(_05327_));
 sky130_fd_sc_hd__clkbuf_1 _25261_ (.A(_05327_),
    .X(_00171_));
 sky130_fd_sc_hd__clkbuf_2 _25262_ (.A(_05224_),
    .X(_05328_));
 sky130_fd_sc_hd__mux2_1 _25263_ (.A0(_05328_),
    .A1(\cpuregs[3][26] ),
    .S(_05324_),
    .X(_05329_));
 sky130_fd_sc_hd__clkbuf_1 _25264_ (.A(_05329_),
    .X(_00172_));
 sky130_fd_sc_hd__clkbuf_2 _25265_ (.A(_05231_),
    .X(_05330_));
 sky130_fd_sc_hd__mux2_1 _25266_ (.A0(_05330_),
    .A1(\cpuregs[3][27] ),
    .S(_05324_),
    .X(_05331_));
 sky130_fd_sc_hd__clkbuf_1 _25267_ (.A(_05331_),
    .X(_00173_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _25268_ (.A(_05239_),
    .X(_05332_));
 sky130_fd_sc_hd__mux2_1 _25269_ (.A0(_05332_),
    .A1(\cpuregs[3][28] ),
    .S(_05324_),
    .X(_05333_));
 sky130_fd_sc_hd__clkbuf_1 _25270_ (.A(_05333_),
    .X(_00174_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _25271_ (.A(_05247_),
    .X(_05334_));
 sky130_fd_sc_hd__mux2_1 _25272_ (.A0(_05334_),
    .A1(\cpuregs[3][29] ),
    .S(_05324_),
    .X(_05335_));
 sky130_fd_sc_hd__clkbuf_1 _25273_ (.A(_05335_),
    .X(_00175_));
 sky130_fd_sc_hd__buf_1 _25274_ (.A(_05255_),
    .X(_05336_));
 sky130_fd_sc_hd__mux2_1 _25275_ (.A0(_05336_),
    .A1(\cpuregs[3][30] ),
    .S(_05271_),
    .X(_05337_));
 sky130_fd_sc_hd__clkbuf_1 _25276_ (.A(_05337_),
    .X(_00176_));
 sky130_fd_sc_hd__buf_1 _25277_ (.A(_05262_),
    .X(_05338_));
 sky130_fd_sc_hd__mux2_1 _25278_ (.A0(_05338_),
    .A1(\cpuregs[3][31] ),
    .S(_05271_),
    .X(_05339_));
 sky130_fd_sc_hd__clkbuf_1 _25279_ (.A(_05339_),
    .X(_00177_));
 sky130_fd_sc_hd__or3_2 _25280_ (.A(\latched_rd[1] ),
    .B(_05267_),
    .C(_04989_),
    .X(_05340_));
 sky130_fd_sc_hd__nor2_1 _25281_ (.A(_04991_),
    .B(_05340_),
    .Y(_05341_));
 sky130_fd_sc_hd__clkbuf_4 _25282_ (.A(_05341_),
    .X(_05342_));
 sky130_fd_sc_hd__buf_2 _25283_ (.A(_05342_),
    .X(_05343_));
 sky130_fd_sc_hd__mux2_1 _25284_ (.A0(\cpuregs[5][0] ),
    .A1(_04988_),
    .S(_05343_),
    .X(_05344_));
 sky130_fd_sc_hd__clkbuf_1 _25285_ (.A(_05344_),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _25286_ (.A0(\cpuregs[5][1] ),
    .A1(_05006_),
    .S(_05343_),
    .X(_05345_));
 sky130_fd_sc_hd__clkbuf_1 _25287_ (.A(_05345_),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _25288_ (.A0(\cpuregs[5][2] ),
    .A1(_05016_),
    .S(_05343_),
    .X(_05346_));
 sky130_fd_sc_hd__clkbuf_1 _25289_ (.A(_05346_),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _25290_ (.A0(\cpuregs[5][3] ),
    .A1(_05023_),
    .S(_05343_),
    .X(_05347_));
 sky130_fd_sc_hd__clkbuf_1 _25291_ (.A(_05347_),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _25292_ (.A0(\cpuregs[5][4] ),
    .A1(_05032_),
    .S(_05343_),
    .X(_05348_));
 sky130_fd_sc_hd__clkbuf_1 _25293_ (.A(_05348_),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _25294_ (.A0(\cpuregs[5][5] ),
    .A1(_05041_),
    .S(_05343_),
    .X(_05349_));
 sky130_fd_sc_hd__clkbuf_1 _25295_ (.A(_05349_),
    .X(_00183_));
 sky130_fd_sc_hd__buf_2 _25296_ (.A(_05342_),
    .X(_05350_));
 sky130_fd_sc_hd__mux2_1 _25297_ (.A0(\cpuregs[5][6] ),
    .A1(_05049_),
    .S(_05350_),
    .X(_05351_));
 sky130_fd_sc_hd__clkbuf_1 _25298_ (.A(_05351_),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _25299_ (.A0(\cpuregs[5][7] ),
    .A1(_05060_),
    .S(_05350_),
    .X(_05352_));
 sky130_fd_sc_hd__clkbuf_1 _25300_ (.A(_05352_),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _25301_ (.A0(\cpuregs[5][8] ),
    .A1(_05069_),
    .S(_05350_),
    .X(_05353_));
 sky130_fd_sc_hd__clkbuf_1 _25302_ (.A(_05353_),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _25303_ (.A0(\cpuregs[5][9] ),
    .A1(_05076_),
    .S(_05350_),
    .X(_05354_));
 sky130_fd_sc_hd__clkbuf_1 _25304_ (.A(_05354_),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _25305_ (.A0(\cpuregs[5][10] ),
    .A1(_05085_),
    .S(_05350_),
    .X(_05355_));
 sky130_fd_sc_hd__clkbuf_1 _25306_ (.A(_05355_),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _25307_ (.A0(\cpuregs[5][11] ),
    .A1(_05095_),
    .S(_05350_),
    .X(_05356_));
 sky130_fd_sc_hd__clkbuf_1 _25308_ (.A(_05356_),
    .X(_00189_));
 sky130_fd_sc_hd__buf_2 _25309_ (.A(_05342_),
    .X(_05357_));
 sky130_fd_sc_hd__mux2_1 _25310_ (.A0(\cpuregs[5][12] ),
    .A1(_05102_),
    .S(_05357_),
    .X(_05358_));
 sky130_fd_sc_hd__clkbuf_1 _25311_ (.A(_05358_),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _25312_ (.A0(\cpuregs[5][13] ),
    .A1(_05113_),
    .S(_05357_),
    .X(_05359_));
 sky130_fd_sc_hd__clkbuf_1 _25313_ (.A(_05359_),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _25314_ (.A0(\cpuregs[5][14] ),
    .A1(_05121_),
    .S(_05357_),
    .X(_05360_));
 sky130_fd_sc_hd__clkbuf_1 _25315_ (.A(_05360_),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _25316_ (.A0(\cpuregs[5][15] ),
    .A1(_05129_),
    .S(_05357_),
    .X(_05361_));
 sky130_fd_sc_hd__clkbuf_1 _25317_ (.A(_05361_),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _25318_ (.A0(\cpuregs[5][16] ),
    .A1(_05138_),
    .S(_05357_),
    .X(_05362_));
 sky130_fd_sc_hd__clkbuf_1 _25319_ (.A(_05362_),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _25320_ (.A0(\cpuregs[5][17] ),
    .A1(_05146_),
    .S(_05357_),
    .X(_05363_));
 sky130_fd_sc_hd__clkbuf_1 _25321_ (.A(_05363_),
    .X(_00195_));
 sky130_fd_sc_hd__buf_2 _25322_ (.A(_05342_),
    .X(_05364_));
 sky130_fd_sc_hd__mux2_1 _25323_ (.A0(\cpuregs[5][18] ),
    .A1(_05154_),
    .S(_05364_),
    .X(_05365_));
 sky130_fd_sc_hd__clkbuf_1 _25324_ (.A(_05365_),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _25325_ (.A0(\cpuregs[5][19] ),
    .A1(_05165_),
    .S(_05364_),
    .X(_05366_));
 sky130_fd_sc_hd__clkbuf_1 _25326_ (.A(_05366_),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _25327_ (.A0(\cpuregs[5][20] ),
    .A1(_05173_),
    .S(_05364_),
    .X(_05367_));
 sky130_fd_sc_hd__clkbuf_1 _25328_ (.A(_05367_),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _25329_ (.A0(\cpuregs[5][21] ),
    .A1(_05182_),
    .S(_05364_),
    .X(_05368_));
 sky130_fd_sc_hd__clkbuf_1 _25330_ (.A(_05368_),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _25331_ (.A0(\cpuregs[5][22] ),
    .A1(_05191_),
    .S(_05364_),
    .X(_05369_));
 sky130_fd_sc_hd__clkbuf_1 _25332_ (.A(_05369_),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _25333_ (.A0(\cpuregs[5][23] ),
    .A1(_05199_),
    .S(_05364_),
    .X(_05370_));
 sky130_fd_sc_hd__clkbuf_1 _25334_ (.A(_05370_),
    .X(_00201_));
 sky130_fd_sc_hd__buf_2 _25335_ (.A(_05341_),
    .X(_05371_));
 sky130_fd_sc_hd__mux2_1 _25336_ (.A0(\cpuregs[5][24] ),
    .A1(_05206_),
    .S(_05371_),
    .X(_05372_));
 sky130_fd_sc_hd__clkbuf_1 _25337_ (.A(_05372_),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _25338_ (.A0(\cpuregs[5][25] ),
    .A1(_05217_),
    .S(_05371_),
    .X(_05373_));
 sky130_fd_sc_hd__clkbuf_1 _25339_ (.A(_05373_),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _25340_ (.A0(\cpuregs[5][26] ),
    .A1(_05225_),
    .S(_05371_),
    .X(_05374_));
 sky130_fd_sc_hd__clkbuf_1 _25341_ (.A(_05374_),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _25342_ (.A0(\cpuregs[5][27] ),
    .A1(_05232_),
    .S(_05371_),
    .X(_05375_));
 sky130_fd_sc_hd__clkbuf_1 _25343_ (.A(_05375_),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _25344_ (.A0(\cpuregs[5][28] ),
    .A1(_05240_),
    .S(_05371_),
    .X(_05376_));
 sky130_fd_sc_hd__clkbuf_1 _25345_ (.A(_05376_),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _25346_ (.A0(\cpuregs[5][29] ),
    .A1(_05248_),
    .S(_05371_),
    .X(_05377_));
 sky130_fd_sc_hd__clkbuf_1 _25347_ (.A(_05377_),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _25348_ (.A0(\cpuregs[5][30] ),
    .A1(_05256_),
    .S(_05342_),
    .X(_05378_));
 sky130_fd_sc_hd__clkbuf_1 _25349_ (.A(_05378_),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _25350_ (.A0(\cpuregs[5][31] ),
    .A1(_05263_),
    .S(_05342_),
    .X(_05379_));
 sky130_fd_sc_hd__clkbuf_1 _25351_ (.A(_05379_),
    .X(_00209_));
 sky130_fd_sc_hd__or3b_1 _25352_ (.A(\latched_rd[0] ),
    .B(_04989_),
    .C_N(\latched_rd[1] ),
    .X(_05380_));
 sky130_fd_sc_hd__clkbuf_2 _25353_ (.A(_05380_),
    .X(_05381_));
 sky130_fd_sc_hd__nor2_1 _25354_ (.A(_04991_),
    .B(_05381_),
    .Y(_05382_));
 sky130_fd_sc_hd__buf_4 _25355_ (.A(_05382_),
    .X(_05383_));
 sky130_fd_sc_hd__buf_2 _25356_ (.A(_05383_),
    .X(_05384_));
 sky130_fd_sc_hd__mux2_1 _25357_ (.A0(\cpuregs[6][0] ),
    .A1(_04988_),
    .S(_05384_),
    .X(_05385_));
 sky130_fd_sc_hd__clkbuf_1 _25358_ (.A(_05385_),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _25359_ (.A0(\cpuregs[6][1] ),
    .A1(_05006_),
    .S(_05384_),
    .X(_05386_));
 sky130_fd_sc_hd__clkbuf_1 _25360_ (.A(_05386_),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _25361_ (.A0(\cpuregs[6][2] ),
    .A1(_05016_),
    .S(_05384_),
    .X(_05387_));
 sky130_fd_sc_hd__clkbuf_1 _25362_ (.A(_05387_),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _25363_ (.A0(\cpuregs[6][3] ),
    .A1(_05023_),
    .S(_05384_),
    .X(_05388_));
 sky130_fd_sc_hd__clkbuf_1 _25364_ (.A(_05388_),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _25365_ (.A0(\cpuregs[6][4] ),
    .A1(_05032_),
    .S(_05384_),
    .X(_05389_));
 sky130_fd_sc_hd__clkbuf_1 _25366_ (.A(_05389_),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _25367_ (.A0(\cpuregs[6][5] ),
    .A1(_05041_),
    .S(_05384_),
    .X(_05390_));
 sky130_fd_sc_hd__clkbuf_1 _25368_ (.A(_05390_),
    .X(_00215_));
 sky130_fd_sc_hd__clkbuf_4 _25369_ (.A(_05383_),
    .X(_05391_));
 sky130_fd_sc_hd__mux2_1 _25370_ (.A0(\cpuregs[6][6] ),
    .A1(_05049_),
    .S(_05391_),
    .X(_05392_));
 sky130_fd_sc_hd__clkbuf_1 _25371_ (.A(_05392_),
    .X(_00216_));
 sky130_fd_sc_hd__mux2_1 _25372_ (.A0(\cpuregs[6][7] ),
    .A1(_05060_),
    .S(_05391_),
    .X(_05393_));
 sky130_fd_sc_hd__clkbuf_1 _25373_ (.A(_05393_),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _25374_ (.A0(\cpuregs[6][8] ),
    .A1(_05069_),
    .S(_05391_),
    .X(_05394_));
 sky130_fd_sc_hd__clkbuf_1 _25375_ (.A(_05394_),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _25376_ (.A0(\cpuregs[6][9] ),
    .A1(_05076_),
    .S(_05391_),
    .X(_05395_));
 sky130_fd_sc_hd__clkbuf_1 _25377_ (.A(_05395_),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_1 _25378_ (.A0(\cpuregs[6][10] ),
    .A1(_05085_),
    .S(_05391_),
    .X(_05396_));
 sky130_fd_sc_hd__clkbuf_1 _25379_ (.A(_05396_),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _25380_ (.A0(\cpuregs[6][11] ),
    .A1(_05095_),
    .S(_05391_),
    .X(_05397_));
 sky130_fd_sc_hd__clkbuf_1 _25381_ (.A(_05397_),
    .X(_00221_));
 sky130_fd_sc_hd__buf_2 _25382_ (.A(_05383_),
    .X(_05398_));
 sky130_fd_sc_hd__mux2_1 _25383_ (.A0(\cpuregs[6][12] ),
    .A1(_05102_),
    .S(_05398_),
    .X(_05399_));
 sky130_fd_sc_hd__clkbuf_1 _25384_ (.A(_05399_),
    .X(_00222_));
 sky130_fd_sc_hd__mux2_1 _25385_ (.A0(\cpuregs[6][13] ),
    .A1(_05113_),
    .S(_05398_),
    .X(_05400_));
 sky130_fd_sc_hd__clkbuf_1 _25386_ (.A(_05400_),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _25387_ (.A0(\cpuregs[6][14] ),
    .A1(_05121_),
    .S(_05398_),
    .X(_05401_));
 sky130_fd_sc_hd__clkbuf_1 _25388_ (.A(_05401_),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_1 _25389_ (.A0(\cpuregs[6][15] ),
    .A1(_05129_),
    .S(_05398_),
    .X(_05402_));
 sky130_fd_sc_hd__clkbuf_1 _25390_ (.A(_05402_),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _25391_ (.A0(\cpuregs[6][16] ),
    .A1(_05138_),
    .S(_05398_),
    .X(_05403_));
 sky130_fd_sc_hd__clkbuf_1 _25392_ (.A(_05403_),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _25393_ (.A0(\cpuregs[6][17] ),
    .A1(_05146_),
    .S(_05398_),
    .X(_05404_));
 sky130_fd_sc_hd__clkbuf_1 _25394_ (.A(_05404_),
    .X(_00227_));
 sky130_fd_sc_hd__buf_2 _25395_ (.A(_05383_),
    .X(_05405_));
 sky130_fd_sc_hd__mux2_1 _25396_ (.A0(\cpuregs[6][18] ),
    .A1(_05154_),
    .S(_05405_),
    .X(_05406_));
 sky130_fd_sc_hd__clkbuf_1 _25397_ (.A(_05406_),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _25398_ (.A0(\cpuregs[6][19] ),
    .A1(_05165_),
    .S(_05405_),
    .X(_05407_));
 sky130_fd_sc_hd__clkbuf_1 _25399_ (.A(_05407_),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _25400_ (.A0(\cpuregs[6][20] ),
    .A1(_05173_),
    .S(_05405_),
    .X(_05408_));
 sky130_fd_sc_hd__clkbuf_1 _25401_ (.A(_05408_),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _25402_ (.A0(\cpuregs[6][21] ),
    .A1(_05182_),
    .S(_05405_),
    .X(_05409_));
 sky130_fd_sc_hd__clkbuf_1 _25403_ (.A(_05409_),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _25404_ (.A0(\cpuregs[6][22] ),
    .A1(_05191_),
    .S(_05405_),
    .X(_05410_));
 sky130_fd_sc_hd__clkbuf_1 _25405_ (.A(_05410_),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _25406_ (.A0(\cpuregs[6][23] ),
    .A1(_05199_),
    .S(_05405_),
    .X(_05411_));
 sky130_fd_sc_hd__clkbuf_1 _25407_ (.A(_05411_),
    .X(_00233_));
 sky130_fd_sc_hd__buf_2 _25408_ (.A(_05382_),
    .X(_05412_));
 sky130_fd_sc_hd__mux2_1 _25409_ (.A0(\cpuregs[6][24] ),
    .A1(_05206_),
    .S(_05412_),
    .X(_05413_));
 sky130_fd_sc_hd__clkbuf_1 _25410_ (.A(_05413_),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _25411_ (.A0(\cpuregs[6][25] ),
    .A1(_05217_),
    .S(_05412_),
    .X(_05414_));
 sky130_fd_sc_hd__clkbuf_1 _25412_ (.A(_05414_),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _25413_ (.A0(\cpuregs[6][26] ),
    .A1(_05225_),
    .S(_05412_),
    .X(_05415_));
 sky130_fd_sc_hd__clkbuf_1 _25414_ (.A(_05415_),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_1 _25415_ (.A0(\cpuregs[6][27] ),
    .A1(_05232_),
    .S(_05412_),
    .X(_05416_));
 sky130_fd_sc_hd__clkbuf_1 _25416_ (.A(_05416_),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _25417_ (.A0(\cpuregs[6][28] ),
    .A1(_05240_),
    .S(_05412_),
    .X(_05417_));
 sky130_fd_sc_hd__clkbuf_1 _25418_ (.A(_05417_),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _25419_ (.A0(\cpuregs[6][29] ),
    .A1(_05248_),
    .S(_05412_),
    .X(_05418_));
 sky130_fd_sc_hd__clkbuf_1 _25420_ (.A(_05418_),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _25421_ (.A0(\cpuregs[6][30] ),
    .A1(_05256_),
    .S(_05383_),
    .X(_05419_));
 sky130_fd_sc_hd__clkbuf_1 _25422_ (.A(_05419_),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _25423_ (.A0(\cpuregs[6][31] ),
    .A1(_05263_),
    .S(_05383_),
    .X(_05420_));
 sky130_fd_sc_hd__clkbuf_1 _25424_ (.A(_05420_),
    .X(_00241_));
 sky130_fd_sc_hd__or2_1 _25425_ (.A(\genblk1.pcpi_mul.active[1] ),
    .B(\genblk1.pcpi_mul.active[0] ),
    .X(_05421_));
 sky130_fd_sc_hd__or3_1 _25426_ (.A(_08140_),
    .B(_08141_),
    .C(_08142_),
    .X(_05422_));
 sky130_fd_sc_hd__or3_4 _25427_ (.A(_08139_),
    .B(_05421_),
    .C(_05422_),
    .X(_05423_));
 sky130_fd_sc_hd__clkbuf_4 _25428_ (.A(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__clkbuf_2 _25429_ (.A(_05424_),
    .X(_05425_));
 sky130_fd_sc_hd__nor2_2 _25430_ (.A(_08143_),
    .B(_05421_),
    .Y(_00773_));
 sky130_fd_sc_hd__and4b_1 _25431_ (.A_N(net239),
    .B(net238),
    .C(_00773_),
    .D(_10260_),
    .X(_05426_));
 sky130_fd_sc_hd__a21o_1 _25432_ (.A1(_13805_),
    .A2(_05425_),
    .B1(_05426_),
    .X(_00242_));
 sky130_fd_sc_hd__nand2_1 _25433_ (.A(net239),
    .B(net238),
    .Y(_05427_));
 sky130_fd_sc_hd__and4_1 _25434_ (.A(_10259_),
    .B(\genblk1.pcpi_mul.instr_any_mulh ),
    .C(_00773_),
    .D(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__a21o_1 _25435_ (.A1(_14565_),
    .A2(_05425_),
    .B1(_05428_),
    .X(_00243_));
 sky130_fd_sc_hd__or2_1 _25436_ (.A(_04991_),
    .B(_05268_),
    .X(_05429_));
 sky130_fd_sc_hd__buf_4 _25437_ (.A(_05429_),
    .X(_05430_));
 sky130_fd_sc_hd__buf_2 _25438_ (.A(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__mux2_1 _25439_ (.A0(_05265_),
    .A1(\cpuregs[7][0] ),
    .S(_05431_),
    .X(_05432_));
 sky130_fd_sc_hd__clkbuf_1 _25440_ (.A(_05432_),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _25441_ (.A0(_05274_),
    .A1(\cpuregs[7][1] ),
    .S(_05431_),
    .X(_05433_));
 sky130_fd_sc_hd__clkbuf_1 _25442_ (.A(_05433_),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _25443_ (.A0(_05276_),
    .A1(\cpuregs[7][2] ),
    .S(_05431_),
    .X(_05434_));
 sky130_fd_sc_hd__clkbuf_1 _25444_ (.A(_05434_),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _25445_ (.A0(_05278_),
    .A1(\cpuregs[7][3] ),
    .S(_05431_),
    .X(_05435_));
 sky130_fd_sc_hd__clkbuf_1 _25446_ (.A(_05435_),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _25447_ (.A0(_05280_),
    .A1(\cpuregs[7][4] ),
    .S(_05431_),
    .X(_05436_));
 sky130_fd_sc_hd__clkbuf_1 _25448_ (.A(_05436_),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _25449_ (.A0(_05282_),
    .A1(\cpuregs[7][5] ),
    .S(_05431_),
    .X(_05437_));
 sky130_fd_sc_hd__clkbuf_1 _25450_ (.A(_05437_),
    .X(_00249_));
 sky130_fd_sc_hd__clkbuf_4 _25451_ (.A(_05430_),
    .X(_05438_));
 sky130_fd_sc_hd__mux2_1 _25452_ (.A0(_05284_),
    .A1(\cpuregs[7][6] ),
    .S(_05438_),
    .X(_05439_));
 sky130_fd_sc_hd__clkbuf_1 _25453_ (.A(_05439_),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _25454_ (.A0(_05287_),
    .A1(\cpuregs[7][7] ),
    .S(_05438_),
    .X(_05440_));
 sky130_fd_sc_hd__clkbuf_1 _25455_ (.A(_05440_),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _25456_ (.A0(_05289_),
    .A1(\cpuregs[7][8] ),
    .S(_05438_),
    .X(_05441_));
 sky130_fd_sc_hd__clkbuf_1 _25457_ (.A(_05441_),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _25458_ (.A0(_05291_),
    .A1(\cpuregs[7][9] ),
    .S(_05438_),
    .X(_05442_));
 sky130_fd_sc_hd__clkbuf_1 _25459_ (.A(_05442_),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _25460_ (.A0(_05293_),
    .A1(\cpuregs[7][10] ),
    .S(_05438_),
    .X(_05443_));
 sky130_fd_sc_hd__clkbuf_1 _25461_ (.A(_05443_),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _25462_ (.A0(_05295_),
    .A1(\cpuregs[7][11] ),
    .S(_05438_),
    .X(_05444_));
 sky130_fd_sc_hd__clkbuf_1 _25463_ (.A(_05444_),
    .X(_00255_));
 sky130_fd_sc_hd__buf_2 _25464_ (.A(_05430_),
    .X(_05445_));
 sky130_fd_sc_hd__mux2_1 _25465_ (.A0(_05297_),
    .A1(\cpuregs[7][12] ),
    .S(_05445_),
    .X(_05446_));
 sky130_fd_sc_hd__clkbuf_1 _25466_ (.A(_05446_),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _25467_ (.A0(_05300_),
    .A1(\cpuregs[7][13] ),
    .S(_05445_),
    .X(_05447_));
 sky130_fd_sc_hd__clkbuf_1 _25468_ (.A(_05447_),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _25469_ (.A0(_05302_),
    .A1(\cpuregs[7][14] ),
    .S(_05445_),
    .X(_05448_));
 sky130_fd_sc_hd__clkbuf_1 _25470_ (.A(_05448_),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _25471_ (.A0(_05304_),
    .A1(\cpuregs[7][15] ),
    .S(_05445_),
    .X(_05449_));
 sky130_fd_sc_hd__clkbuf_1 _25472_ (.A(_05449_),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _25473_ (.A0(_05306_),
    .A1(\cpuregs[7][16] ),
    .S(_05445_),
    .X(_05450_));
 sky130_fd_sc_hd__clkbuf_1 _25474_ (.A(_05450_),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _25475_ (.A0(_05308_),
    .A1(\cpuregs[7][17] ),
    .S(_05445_),
    .X(_05451_));
 sky130_fd_sc_hd__clkbuf_1 _25476_ (.A(_05451_),
    .X(_00261_));
 sky130_fd_sc_hd__buf_2 _25477_ (.A(_05430_),
    .X(_05452_));
 sky130_fd_sc_hd__mux2_1 _25478_ (.A0(_05310_),
    .A1(\cpuregs[7][18] ),
    .S(_05452_),
    .X(_05453_));
 sky130_fd_sc_hd__clkbuf_1 _25479_ (.A(_05453_),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _25480_ (.A0(_05313_),
    .A1(\cpuregs[7][19] ),
    .S(_05452_),
    .X(_05454_));
 sky130_fd_sc_hd__clkbuf_1 _25481_ (.A(_05454_),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _25482_ (.A0(_05315_),
    .A1(\cpuregs[7][20] ),
    .S(_05452_),
    .X(_05455_));
 sky130_fd_sc_hd__clkbuf_1 _25483_ (.A(_05455_),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _25484_ (.A0(_05317_),
    .A1(\cpuregs[7][21] ),
    .S(_05452_),
    .X(_05456_));
 sky130_fd_sc_hd__clkbuf_1 _25485_ (.A(_05456_),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _25486_ (.A0(_05319_),
    .A1(\cpuregs[7][22] ),
    .S(_05452_),
    .X(_05457_));
 sky130_fd_sc_hd__clkbuf_1 _25487_ (.A(_05457_),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _25488_ (.A0(_05321_),
    .A1(\cpuregs[7][23] ),
    .S(_05452_),
    .X(_05458_));
 sky130_fd_sc_hd__clkbuf_1 _25489_ (.A(_05458_),
    .X(_00267_));
 sky130_fd_sc_hd__buf_2 _25490_ (.A(_05429_),
    .X(_05459_));
 sky130_fd_sc_hd__mux2_1 _25491_ (.A0(_05323_),
    .A1(\cpuregs[7][24] ),
    .S(_05459_),
    .X(_05460_));
 sky130_fd_sc_hd__clkbuf_1 _25492_ (.A(_05460_),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _25493_ (.A0(_05326_),
    .A1(\cpuregs[7][25] ),
    .S(_05459_),
    .X(_05461_));
 sky130_fd_sc_hd__clkbuf_1 _25494_ (.A(_05461_),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _25495_ (.A0(_05328_),
    .A1(\cpuregs[7][26] ),
    .S(_05459_),
    .X(_05462_));
 sky130_fd_sc_hd__clkbuf_1 _25496_ (.A(_05462_),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _25497_ (.A0(_05330_),
    .A1(\cpuregs[7][27] ),
    .S(_05459_),
    .X(_05463_));
 sky130_fd_sc_hd__clkbuf_1 _25498_ (.A(_05463_),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _25499_ (.A0(_05332_),
    .A1(\cpuregs[7][28] ),
    .S(_05459_),
    .X(_05464_));
 sky130_fd_sc_hd__clkbuf_1 _25500_ (.A(_05464_),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _25501_ (.A0(_05334_),
    .A1(\cpuregs[7][29] ),
    .S(_05459_),
    .X(_05465_));
 sky130_fd_sc_hd__clkbuf_1 _25502_ (.A(_05465_),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _25503_ (.A0(_05336_),
    .A1(\cpuregs[7][30] ),
    .S(_05430_),
    .X(_05466_));
 sky130_fd_sc_hd__clkbuf_1 _25504_ (.A(_05466_),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _25505_ (.A0(_05338_),
    .A1(\cpuregs[7][31] ),
    .S(_05430_),
    .X(_05467_));
 sky130_fd_sc_hd__clkbuf_1 _25506_ (.A(_05467_),
    .X(_00275_));
 sky130_fd_sc_hd__or3b_1 _25507_ (.A(\latched_rd[2] ),
    .B(\latched_rd[4] ),
    .C_N(\latched_rd[3] ),
    .X(_05468_));
 sky130_fd_sc_hd__nor2_1 _25508_ (.A(_04990_),
    .B(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__clkbuf_4 _25509_ (.A(_05469_),
    .X(_05470_));
 sky130_fd_sc_hd__buf_2 _25510_ (.A(_05470_),
    .X(_05471_));
 sky130_fd_sc_hd__mux2_1 _25511_ (.A0(\cpuregs[8][0] ),
    .A1(_04988_),
    .S(_05471_),
    .X(_05472_));
 sky130_fd_sc_hd__clkbuf_1 _25512_ (.A(_05472_),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _25513_ (.A0(\cpuregs[8][1] ),
    .A1(_05006_),
    .S(_05471_),
    .X(_05473_));
 sky130_fd_sc_hd__clkbuf_1 _25514_ (.A(_05473_),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _25515_ (.A0(\cpuregs[8][2] ),
    .A1(_05016_),
    .S(_05471_),
    .X(_05474_));
 sky130_fd_sc_hd__clkbuf_1 _25516_ (.A(_05474_),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _25517_ (.A0(\cpuregs[8][3] ),
    .A1(_05023_),
    .S(_05471_),
    .X(_05475_));
 sky130_fd_sc_hd__clkbuf_1 _25518_ (.A(_05475_),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _25519_ (.A0(\cpuregs[8][4] ),
    .A1(_05032_),
    .S(_05471_),
    .X(_05476_));
 sky130_fd_sc_hd__clkbuf_1 _25520_ (.A(_05476_),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _25521_ (.A0(\cpuregs[8][5] ),
    .A1(_05041_),
    .S(_05471_),
    .X(_05477_));
 sky130_fd_sc_hd__clkbuf_1 _25522_ (.A(_05477_),
    .X(_00281_));
 sky130_fd_sc_hd__clkbuf_4 _25523_ (.A(_05470_),
    .X(_05478_));
 sky130_fd_sc_hd__mux2_1 _25524_ (.A0(\cpuregs[8][6] ),
    .A1(_05049_),
    .S(_05478_),
    .X(_05479_));
 sky130_fd_sc_hd__clkbuf_1 _25525_ (.A(_05479_),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _25526_ (.A0(\cpuregs[8][7] ),
    .A1(_05060_),
    .S(_05478_),
    .X(_05480_));
 sky130_fd_sc_hd__clkbuf_1 _25527_ (.A(_05480_),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _25528_ (.A0(\cpuregs[8][8] ),
    .A1(_05069_),
    .S(_05478_),
    .X(_05481_));
 sky130_fd_sc_hd__clkbuf_1 _25529_ (.A(_05481_),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _25530_ (.A0(\cpuregs[8][9] ),
    .A1(_05076_),
    .S(_05478_),
    .X(_05482_));
 sky130_fd_sc_hd__clkbuf_1 _25531_ (.A(_05482_),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _25532_ (.A0(\cpuregs[8][10] ),
    .A1(_05085_),
    .S(_05478_),
    .X(_05483_));
 sky130_fd_sc_hd__clkbuf_1 _25533_ (.A(_05483_),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _25534_ (.A0(\cpuregs[8][11] ),
    .A1(_05095_),
    .S(_05478_),
    .X(_05484_));
 sky130_fd_sc_hd__clkbuf_1 _25535_ (.A(_05484_),
    .X(_00287_));
 sky130_fd_sc_hd__clkbuf_4 _25536_ (.A(_05470_),
    .X(_05485_));
 sky130_fd_sc_hd__mux2_1 _25537_ (.A0(\cpuregs[8][12] ),
    .A1(_05102_),
    .S(_05485_),
    .X(_05486_));
 sky130_fd_sc_hd__clkbuf_1 _25538_ (.A(_05486_),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _25539_ (.A0(\cpuregs[8][13] ),
    .A1(_05113_),
    .S(_05485_),
    .X(_05487_));
 sky130_fd_sc_hd__clkbuf_1 _25540_ (.A(_05487_),
    .X(_00289_));
 sky130_fd_sc_hd__mux2_1 _25541_ (.A0(\cpuregs[8][14] ),
    .A1(_05121_),
    .S(_05485_),
    .X(_05488_));
 sky130_fd_sc_hd__clkbuf_1 _25542_ (.A(_05488_),
    .X(_00290_));
 sky130_fd_sc_hd__mux2_1 _25543_ (.A0(\cpuregs[8][15] ),
    .A1(_05129_),
    .S(_05485_),
    .X(_05489_));
 sky130_fd_sc_hd__clkbuf_1 _25544_ (.A(_05489_),
    .X(_00291_));
 sky130_fd_sc_hd__mux2_1 _25545_ (.A0(\cpuregs[8][16] ),
    .A1(_05138_),
    .S(_05485_),
    .X(_05490_));
 sky130_fd_sc_hd__clkbuf_1 _25546_ (.A(_05490_),
    .X(_00292_));
 sky130_fd_sc_hd__mux2_1 _25547_ (.A0(\cpuregs[8][17] ),
    .A1(_05146_),
    .S(_05485_),
    .X(_05491_));
 sky130_fd_sc_hd__clkbuf_1 _25548_ (.A(_05491_),
    .X(_00293_));
 sky130_fd_sc_hd__buf_2 _25549_ (.A(_05470_),
    .X(_05492_));
 sky130_fd_sc_hd__mux2_1 _25550_ (.A0(\cpuregs[8][18] ),
    .A1(_05154_),
    .S(_05492_),
    .X(_05493_));
 sky130_fd_sc_hd__clkbuf_1 _25551_ (.A(_05493_),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _25552_ (.A0(\cpuregs[8][19] ),
    .A1(_05165_),
    .S(_05492_),
    .X(_05494_));
 sky130_fd_sc_hd__clkbuf_1 _25553_ (.A(_05494_),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_1 _25554_ (.A0(\cpuregs[8][20] ),
    .A1(_05173_),
    .S(_05492_),
    .X(_05495_));
 sky130_fd_sc_hd__clkbuf_1 _25555_ (.A(_05495_),
    .X(_00296_));
 sky130_fd_sc_hd__mux2_1 _25556_ (.A0(\cpuregs[8][21] ),
    .A1(_05182_),
    .S(_05492_),
    .X(_05496_));
 sky130_fd_sc_hd__clkbuf_1 _25557_ (.A(_05496_),
    .X(_00297_));
 sky130_fd_sc_hd__mux2_1 _25558_ (.A0(\cpuregs[8][22] ),
    .A1(_05191_),
    .S(_05492_),
    .X(_05497_));
 sky130_fd_sc_hd__clkbuf_1 _25559_ (.A(_05497_),
    .X(_00298_));
 sky130_fd_sc_hd__mux2_1 _25560_ (.A0(\cpuregs[8][23] ),
    .A1(_05199_),
    .S(_05492_),
    .X(_05498_));
 sky130_fd_sc_hd__clkbuf_1 _25561_ (.A(_05498_),
    .X(_00299_));
 sky130_fd_sc_hd__clkbuf_4 _25562_ (.A(_05469_),
    .X(_05499_));
 sky130_fd_sc_hd__mux2_1 _25563_ (.A0(\cpuregs[8][24] ),
    .A1(_05206_),
    .S(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__clkbuf_1 _25564_ (.A(_05500_),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _25565_ (.A0(\cpuregs[8][25] ),
    .A1(_05217_),
    .S(_05499_),
    .X(_05501_));
 sky130_fd_sc_hd__clkbuf_1 _25566_ (.A(_05501_),
    .X(_00301_));
 sky130_fd_sc_hd__mux2_1 _25567_ (.A0(\cpuregs[8][26] ),
    .A1(_05225_),
    .S(_05499_),
    .X(_05502_));
 sky130_fd_sc_hd__clkbuf_1 _25568_ (.A(_05502_),
    .X(_00302_));
 sky130_fd_sc_hd__mux2_1 _25569_ (.A0(\cpuregs[8][27] ),
    .A1(_05232_),
    .S(_05499_),
    .X(_05503_));
 sky130_fd_sc_hd__clkbuf_1 _25570_ (.A(_05503_),
    .X(_00303_));
 sky130_fd_sc_hd__mux2_1 _25571_ (.A0(\cpuregs[8][28] ),
    .A1(_05240_),
    .S(_05499_),
    .X(_05504_));
 sky130_fd_sc_hd__clkbuf_1 _25572_ (.A(_05504_),
    .X(_00304_));
 sky130_fd_sc_hd__mux2_1 _25573_ (.A0(\cpuregs[8][29] ),
    .A1(_05248_),
    .S(_05499_),
    .X(_05505_));
 sky130_fd_sc_hd__clkbuf_1 _25574_ (.A(_05505_),
    .X(_00305_));
 sky130_fd_sc_hd__mux2_1 _25575_ (.A0(\cpuregs[8][30] ),
    .A1(_05256_),
    .S(_05470_),
    .X(_05506_));
 sky130_fd_sc_hd__clkbuf_1 _25576_ (.A(_05506_),
    .X(_00306_));
 sky130_fd_sc_hd__mux2_1 _25577_ (.A0(\cpuregs[8][31] ),
    .A1(_05263_),
    .S(_05470_),
    .X(_05507_));
 sky130_fd_sc_hd__clkbuf_1 _25578_ (.A(_05507_),
    .X(_00307_));
 sky130_fd_sc_hd__clkbuf_2 _25579_ (.A(_08155_),
    .X(_05508_));
 sky130_fd_sc_hd__clkbuf_2 _25580_ (.A(_05508_),
    .X(_05509_));
 sky130_fd_sc_hd__clkbuf_2 _25581_ (.A(_05509_),
    .X(_05510_));
 sky130_fd_sc_hd__mux2_1 _25582_ (.A0(net49),
    .A1(\mem_rdata_q[24] ),
    .S(_05510_),
    .X(_05511_));
 sky130_fd_sc_hd__clkbuf_1 _25583_ (.A(_05511_),
    .X(_00637_));
 sky130_fd_sc_hd__and3_1 _25584_ (.A(_08522_),
    .B(_08146_),
    .C(_08157_),
    .X(_05512_));
 sky130_fd_sc_hd__buf_2 _25585_ (.A(_05512_),
    .X(_05513_));
 sky130_fd_sc_hd__mux2_1 _25586_ (.A0(\decoded_imm_uj[4] ),
    .A1(_00637_),
    .S(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__clkbuf_1 _25587_ (.A(_05514_),
    .X(_00308_));
 sky130_fd_sc_hd__mux2_1 _25588_ (.A0(net50),
    .A1(\mem_rdata_q[25] ),
    .S(_08155_),
    .X(_05515_));
 sky130_fd_sc_hd__buf_1 _25589_ (.A(_05515_),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_1 _25590_ (.A0(\decoded_imm_uj[5] ),
    .A1(_00638_),
    .S(_05513_),
    .X(_05516_));
 sky130_fd_sc_hd__clkbuf_1 _25591_ (.A(_05516_),
    .X(_00309_));
 sky130_fd_sc_hd__mux2_1 _25592_ (.A0(net51),
    .A1(\mem_rdata_q[26] ),
    .S(_05509_),
    .X(_05517_));
 sky130_fd_sc_hd__buf_1 _25593_ (.A(_05517_),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _25594_ (.A0(\decoded_imm_uj[6] ),
    .A1(_00639_),
    .S(_05513_),
    .X(_05518_));
 sky130_fd_sc_hd__clkbuf_1 _25595_ (.A(_05518_),
    .X(_00310_));
 sky130_fd_sc_hd__mux2_1 _25596_ (.A0(net52),
    .A1(\mem_rdata_q[27] ),
    .S(_05509_),
    .X(_05519_));
 sky130_fd_sc_hd__buf_1 _25597_ (.A(_05519_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _25598_ (.A0(\decoded_imm_uj[7] ),
    .A1(_00640_),
    .S(_05513_),
    .X(_05520_));
 sky130_fd_sc_hd__clkbuf_1 _25599_ (.A(_05520_),
    .X(_00311_));
 sky130_fd_sc_hd__mux2_1 _25600_ (.A0(net53),
    .A1(\mem_rdata_q[28] ),
    .S(_05509_),
    .X(_05521_));
 sky130_fd_sc_hd__buf_1 _25601_ (.A(_05521_),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_1 _25602_ (.A0(\decoded_imm_uj[8] ),
    .A1(_00641_),
    .S(_05513_),
    .X(_05522_));
 sky130_fd_sc_hd__clkbuf_1 _25603_ (.A(_05522_),
    .X(_00312_));
 sky130_fd_sc_hd__buf_2 _25604_ (.A(_08155_),
    .X(_05523_));
 sky130_fd_sc_hd__mux2_1 _25605_ (.A0(net54),
    .A1(\mem_rdata_q[29] ),
    .S(_05523_),
    .X(_05524_));
 sky130_fd_sc_hd__buf_1 _25606_ (.A(_05524_),
    .X(_00642_));
 sky130_fd_sc_hd__clkbuf_2 _25607_ (.A(_05512_),
    .X(_05525_));
 sky130_fd_sc_hd__mux2_1 _25608_ (.A0(\decoded_imm_uj[9] ),
    .A1(_00642_),
    .S(_05525_),
    .X(_05526_));
 sky130_fd_sc_hd__clkbuf_1 _25609_ (.A(_05526_),
    .X(_00313_));
 sky130_fd_sc_hd__mux2_1 _25610_ (.A0(net56),
    .A1(\mem_rdata_q[30] ),
    .S(_05523_),
    .X(_05527_));
 sky130_fd_sc_hd__buf_1 _25611_ (.A(_05527_),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _25612_ (.A0(\decoded_imm_uj[10] ),
    .A1(_00643_),
    .S(_05525_),
    .X(_05528_));
 sky130_fd_sc_hd__clkbuf_1 _25613_ (.A(_05528_),
    .X(_00314_));
 sky130_fd_sc_hd__buf_2 _25614_ (.A(_05508_),
    .X(_05529_));
 sky130_fd_sc_hd__mux2_1 _25615_ (.A0(net36),
    .A1(\mem_rdata_q[12] ),
    .S(_05529_),
    .X(_05530_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _25616_ (.A(_05530_),
    .X(_00625_));
 sky130_fd_sc_hd__mux2_1 _25617_ (.A0(\decoded_imm_uj[12] ),
    .A1(_00625_),
    .S(_05525_),
    .X(_05531_));
 sky130_fd_sc_hd__clkbuf_1 _25618_ (.A(_05531_),
    .X(_00315_));
 sky130_fd_sc_hd__mux2_1 _25619_ (.A0(net37),
    .A1(\mem_rdata_q[13] ),
    .S(_05529_),
    .X(_05532_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _25620_ (.A(_05532_),
    .X(_00626_));
 sky130_fd_sc_hd__mux2_1 _25621_ (.A0(\decoded_imm_uj[13] ),
    .A1(_00626_),
    .S(_05525_),
    .X(_05533_));
 sky130_fd_sc_hd__clkbuf_1 _25622_ (.A(_05533_),
    .X(_00316_));
 sky130_fd_sc_hd__mux2_1 _25623_ (.A0(net38),
    .A1(\mem_rdata_q[14] ),
    .S(_05529_),
    .X(_05534_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _25624_ (.A(_05534_),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_1 _25625_ (.A0(\decoded_imm_uj[14] ),
    .A1(_00627_),
    .S(_05525_),
    .X(_05535_));
 sky130_fd_sc_hd__clkbuf_1 _25626_ (.A(_05535_),
    .X(_00317_));
 sky130_fd_sc_hd__clkbuf_2 _25627_ (.A(_08536_),
    .X(_05536_));
 sky130_fd_sc_hd__buf_2 _25628_ (.A(_05512_),
    .X(_05537_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _25629_ (.A(_05537_),
    .X(_05538_));
 sky130_fd_sc_hd__mux2_1 _25630_ (.A0(net39),
    .A1(\mem_rdata_q[15] ),
    .S(_05510_),
    .X(_05539_));
 sky130_fd_sc_hd__buf_1 _25631_ (.A(_05539_),
    .X(_00628_));
 sky130_fd_sc_hd__nand2_1 _25632_ (.A(_05538_),
    .B(_00628_),
    .Y(_05540_));
 sky130_fd_sc_hd__a21bo_1 _25633_ (.A1(\decoded_imm_uj[15] ),
    .A2(_05536_),
    .B1_N(_05540_),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _25634_ (.A0(net40),
    .A1(\mem_rdata_q[16] ),
    .S(_05510_),
    .X(_05541_));
 sky130_fd_sc_hd__clkbuf_1 _25635_ (.A(_05541_),
    .X(_00629_));
 sky130_fd_sc_hd__nand2_1 _25636_ (.A(_05538_),
    .B(_00629_),
    .Y(_05542_));
 sky130_fd_sc_hd__a21bo_1 _25637_ (.A1(\decoded_imm_uj[16] ),
    .A2(_05536_),
    .B1_N(_05542_),
    .X(_00319_));
 sky130_fd_sc_hd__mux2_1 _25638_ (.A0(net41),
    .A1(\mem_rdata_q[17] ),
    .S(_05510_),
    .X(_05543_));
 sky130_fd_sc_hd__clkbuf_1 _25639_ (.A(_05543_),
    .X(_00630_));
 sky130_fd_sc_hd__nand2_1 _25640_ (.A(_05538_),
    .B(_00630_),
    .Y(_05544_));
 sky130_fd_sc_hd__a21bo_1 _25641_ (.A1(\decoded_imm_uj[17] ),
    .A2(_05536_),
    .B1_N(_05544_),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _25642_ (.A0(net42),
    .A1(\mem_rdata_q[18] ),
    .S(_05510_),
    .X(_05545_));
 sky130_fd_sc_hd__clkbuf_1 _25643_ (.A(_05545_),
    .X(_00631_));
 sky130_fd_sc_hd__nand2_1 _25644_ (.A(_05538_),
    .B(_00631_),
    .Y(_05546_));
 sky130_fd_sc_hd__a21bo_1 _25645_ (.A1(\decoded_imm_uj[18] ),
    .A2(_05536_),
    .B1_N(_05546_),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _25646_ (.A0(net43),
    .A1(\mem_rdata_q[19] ),
    .S(_05510_),
    .X(_05547_));
 sky130_fd_sc_hd__clkbuf_1 _25647_ (.A(_05547_),
    .X(_00632_));
 sky130_fd_sc_hd__nor2_1 _25648_ (.A(_08536_),
    .B(_00632_),
    .Y(_05548_));
 sky130_fd_sc_hd__o21ba_1 _25649_ (.A1(\decoded_imm_uj[19] ),
    .A2(_05538_),
    .B1_N(_05548_),
    .X(_00322_));
 sky130_fd_sc_hd__buf_2 _25650_ (.A(\decoded_imm_uj[20] ),
    .X(_05549_));
 sky130_fd_sc_hd__clkbuf_2 _25651_ (.A(_05549_),
    .X(_05550_));
 sky130_fd_sc_hd__clkbuf_2 _25652_ (.A(_05550_),
    .X(_05551_));
 sky130_fd_sc_hd__clkbuf_4 _25653_ (.A(_05551_),
    .X(_05552_));
 sky130_fd_sc_hd__mux2_1 _25654_ (.A0(net57),
    .A1(\mem_rdata_q[31] ),
    .S(_05508_),
    .X(_05553_));
 sky130_fd_sc_hd__buf_1 _25655_ (.A(_05553_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _25656_ (.A0(_05552_),
    .A1(_00644_),
    .S(_05525_),
    .X(_05554_));
 sky130_fd_sc_hd__buf_1 _25657_ (.A(_05554_),
    .X(_00323_));
 sky130_fd_sc_hd__clkbuf_1 _25658_ (.A(\cpuregs[0][0] ),
    .X(_05555_));
 sky130_fd_sc_hd__clkbuf_1 _25659_ (.A(_05555_),
    .X(_00324_));
 sky130_fd_sc_hd__clkbuf_1 _25660_ (.A(\cpuregs[0][1] ),
    .X(_05556_));
 sky130_fd_sc_hd__clkbuf_1 _25661_ (.A(_05556_),
    .X(_00325_));
 sky130_fd_sc_hd__clkbuf_1 _25662_ (.A(\cpuregs[0][2] ),
    .X(_05557_));
 sky130_fd_sc_hd__clkbuf_1 _25663_ (.A(_05557_),
    .X(_00326_));
 sky130_fd_sc_hd__clkbuf_1 _25664_ (.A(\cpuregs[0][3] ),
    .X(_05558_));
 sky130_fd_sc_hd__clkbuf_1 _25665_ (.A(_05558_),
    .X(_00327_));
 sky130_fd_sc_hd__clkbuf_1 _25666_ (.A(\cpuregs[0][4] ),
    .X(_05559_));
 sky130_fd_sc_hd__clkbuf_1 _25667_ (.A(_05559_),
    .X(_00328_));
 sky130_fd_sc_hd__clkbuf_1 _25668_ (.A(\cpuregs[0][5] ),
    .X(_05560_));
 sky130_fd_sc_hd__clkbuf_1 _25669_ (.A(_05560_),
    .X(_00329_));
 sky130_fd_sc_hd__clkbuf_1 _25670_ (.A(\cpuregs[0][6] ),
    .X(_05561_));
 sky130_fd_sc_hd__clkbuf_1 _25671_ (.A(_05561_),
    .X(_00330_));
 sky130_fd_sc_hd__clkbuf_1 _25672_ (.A(\cpuregs[0][7] ),
    .X(_05562_));
 sky130_fd_sc_hd__clkbuf_1 _25673_ (.A(_05562_),
    .X(_00331_));
 sky130_fd_sc_hd__clkbuf_1 _25674_ (.A(\cpuregs[0][8] ),
    .X(_05563_));
 sky130_fd_sc_hd__clkbuf_1 _25675_ (.A(_05563_),
    .X(_00332_));
 sky130_fd_sc_hd__clkbuf_1 _25676_ (.A(\cpuregs[0][9] ),
    .X(_05564_));
 sky130_fd_sc_hd__clkbuf_1 _25677_ (.A(_05564_),
    .X(_00333_));
 sky130_fd_sc_hd__clkbuf_1 _25678_ (.A(\cpuregs[0][10] ),
    .X(_05565_));
 sky130_fd_sc_hd__clkbuf_1 _25679_ (.A(_05565_),
    .X(_00334_));
 sky130_fd_sc_hd__clkbuf_1 _25680_ (.A(\cpuregs[0][11] ),
    .X(_05566_));
 sky130_fd_sc_hd__clkbuf_1 _25681_ (.A(_05566_),
    .X(_00335_));
 sky130_fd_sc_hd__clkbuf_1 _25682_ (.A(\cpuregs[0][12] ),
    .X(_05567_));
 sky130_fd_sc_hd__clkbuf_1 _25683_ (.A(_05567_),
    .X(_00336_));
 sky130_fd_sc_hd__clkbuf_1 _25684_ (.A(\cpuregs[0][13] ),
    .X(_05568_));
 sky130_fd_sc_hd__clkbuf_1 _25685_ (.A(_05568_),
    .X(_00337_));
 sky130_fd_sc_hd__clkbuf_1 _25686_ (.A(\cpuregs[0][14] ),
    .X(_05569_));
 sky130_fd_sc_hd__clkbuf_1 _25687_ (.A(_05569_),
    .X(_00338_));
 sky130_fd_sc_hd__clkbuf_1 _25688_ (.A(\cpuregs[0][15] ),
    .X(_05570_));
 sky130_fd_sc_hd__clkbuf_1 _25689_ (.A(_05570_),
    .X(_00339_));
 sky130_fd_sc_hd__clkbuf_1 _25690_ (.A(\cpuregs[0][16] ),
    .X(_05571_));
 sky130_fd_sc_hd__clkbuf_1 _25691_ (.A(_05571_),
    .X(_00340_));
 sky130_fd_sc_hd__clkbuf_1 _25692_ (.A(\cpuregs[0][17] ),
    .X(_05572_));
 sky130_fd_sc_hd__clkbuf_1 _25693_ (.A(_05572_),
    .X(_00341_));
 sky130_fd_sc_hd__clkbuf_1 _25694_ (.A(\cpuregs[0][18] ),
    .X(_05573_));
 sky130_fd_sc_hd__clkbuf_1 _25695_ (.A(_05573_),
    .X(_00342_));
 sky130_fd_sc_hd__clkbuf_1 _25696_ (.A(\cpuregs[0][19] ),
    .X(_05574_));
 sky130_fd_sc_hd__clkbuf_1 _25697_ (.A(_05574_),
    .X(_00343_));
 sky130_fd_sc_hd__clkbuf_1 _25698_ (.A(\cpuregs[0][20] ),
    .X(_05575_));
 sky130_fd_sc_hd__clkbuf_1 _25699_ (.A(_05575_),
    .X(_00344_));
 sky130_fd_sc_hd__clkbuf_1 _25700_ (.A(\cpuregs[0][21] ),
    .X(_05576_));
 sky130_fd_sc_hd__clkbuf_1 _25701_ (.A(_05576_),
    .X(_00345_));
 sky130_fd_sc_hd__clkbuf_1 _25702_ (.A(\cpuregs[0][22] ),
    .X(_05577_));
 sky130_fd_sc_hd__clkbuf_1 _25703_ (.A(_05577_),
    .X(_00346_));
 sky130_fd_sc_hd__clkbuf_1 _25704_ (.A(\cpuregs[0][23] ),
    .X(_05578_));
 sky130_fd_sc_hd__clkbuf_1 _25705_ (.A(_05578_),
    .X(_00347_));
 sky130_fd_sc_hd__clkbuf_1 _25706_ (.A(\cpuregs[0][24] ),
    .X(_05579_));
 sky130_fd_sc_hd__clkbuf_1 _25707_ (.A(_05579_),
    .X(_00348_));
 sky130_fd_sc_hd__clkbuf_1 _25708_ (.A(\cpuregs[0][25] ),
    .X(_05580_));
 sky130_fd_sc_hd__clkbuf_1 _25709_ (.A(_05580_),
    .X(_00349_));
 sky130_fd_sc_hd__clkbuf_1 _25710_ (.A(\cpuregs[0][26] ),
    .X(_05581_));
 sky130_fd_sc_hd__clkbuf_1 _25711_ (.A(_05581_),
    .X(_00350_));
 sky130_fd_sc_hd__clkbuf_1 _25712_ (.A(\cpuregs[0][27] ),
    .X(_05582_));
 sky130_fd_sc_hd__clkbuf_1 _25713_ (.A(_05582_),
    .X(_00351_));
 sky130_fd_sc_hd__clkbuf_1 _25714_ (.A(\cpuregs[0][28] ),
    .X(_05583_));
 sky130_fd_sc_hd__clkbuf_1 _25715_ (.A(_05583_),
    .X(_00352_));
 sky130_fd_sc_hd__clkbuf_1 _25716_ (.A(\cpuregs[0][29] ),
    .X(_05584_));
 sky130_fd_sc_hd__clkbuf_1 _25717_ (.A(_05584_),
    .X(_00353_));
 sky130_fd_sc_hd__clkbuf_1 _25718_ (.A(\cpuregs[0][30] ),
    .X(_05585_));
 sky130_fd_sc_hd__clkbuf_1 _25719_ (.A(_05585_),
    .X(_00354_));
 sky130_fd_sc_hd__clkbuf_1 _25720_ (.A(\cpuregs[0][31] ),
    .X(_05586_));
 sky130_fd_sc_hd__clkbuf_1 _25721_ (.A(_05586_),
    .X(_00355_));
 sky130_fd_sc_hd__nor2_1 _25722_ (.A(_05381_),
    .B(_05468_),
    .Y(_05587_));
 sky130_fd_sc_hd__clkbuf_4 _25723_ (.A(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__buf_2 _25724_ (.A(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__mux2_1 _25725_ (.A0(\cpuregs[10][0] ),
    .A1(_04988_),
    .S(_05589_),
    .X(_05590_));
 sky130_fd_sc_hd__clkbuf_1 _25726_ (.A(_05590_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _25727_ (.A0(\cpuregs[10][1] ),
    .A1(_05006_),
    .S(_05589_),
    .X(_05591_));
 sky130_fd_sc_hd__clkbuf_1 _25728_ (.A(_05591_),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _25729_ (.A0(\cpuregs[10][2] ),
    .A1(_05016_),
    .S(_05589_),
    .X(_05592_));
 sky130_fd_sc_hd__clkbuf_1 _25730_ (.A(_05592_),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_1 _25731_ (.A0(\cpuregs[10][3] ),
    .A1(_05023_),
    .S(_05589_),
    .X(_05593_));
 sky130_fd_sc_hd__clkbuf_1 _25732_ (.A(_05593_),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_1 _25733_ (.A0(\cpuregs[10][4] ),
    .A1(_05032_),
    .S(_05589_),
    .X(_05594_));
 sky130_fd_sc_hd__clkbuf_1 _25734_ (.A(_05594_),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _25735_ (.A0(\cpuregs[10][5] ),
    .A1(_05041_),
    .S(_05589_),
    .X(_05595_));
 sky130_fd_sc_hd__clkbuf_1 _25736_ (.A(_05595_),
    .X(_00361_));
 sky130_fd_sc_hd__buf_2 _25737_ (.A(_05588_),
    .X(_05596_));
 sky130_fd_sc_hd__mux2_1 _25738_ (.A0(\cpuregs[10][6] ),
    .A1(_05049_),
    .S(_05596_),
    .X(_05597_));
 sky130_fd_sc_hd__clkbuf_1 _25739_ (.A(_05597_),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _25740_ (.A0(\cpuregs[10][7] ),
    .A1(_05060_),
    .S(_05596_),
    .X(_05598_));
 sky130_fd_sc_hd__clkbuf_1 _25741_ (.A(_05598_),
    .X(_00363_));
 sky130_fd_sc_hd__mux2_1 _25742_ (.A0(\cpuregs[10][8] ),
    .A1(_05069_),
    .S(_05596_),
    .X(_05599_));
 sky130_fd_sc_hd__clkbuf_1 _25743_ (.A(_05599_),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _25744_ (.A0(\cpuregs[10][9] ),
    .A1(_05076_),
    .S(_05596_),
    .X(_05600_));
 sky130_fd_sc_hd__clkbuf_1 _25745_ (.A(_05600_),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_1 _25746_ (.A0(\cpuregs[10][10] ),
    .A1(_05085_),
    .S(_05596_),
    .X(_05601_));
 sky130_fd_sc_hd__clkbuf_1 _25747_ (.A(_05601_),
    .X(_00366_));
 sky130_fd_sc_hd__mux2_1 _25748_ (.A0(\cpuregs[10][11] ),
    .A1(_05095_),
    .S(_05596_),
    .X(_05602_));
 sky130_fd_sc_hd__clkbuf_1 _25749_ (.A(_05602_),
    .X(_00367_));
 sky130_fd_sc_hd__buf_2 _25750_ (.A(_05588_),
    .X(_05603_));
 sky130_fd_sc_hd__mux2_1 _25751_ (.A0(\cpuregs[10][12] ),
    .A1(_05102_),
    .S(_05603_),
    .X(_05604_));
 sky130_fd_sc_hd__clkbuf_1 _25752_ (.A(_05604_),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _25753_ (.A0(\cpuregs[10][13] ),
    .A1(_05113_),
    .S(_05603_),
    .X(_05605_));
 sky130_fd_sc_hd__clkbuf_1 _25754_ (.A(_05605_),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_1 _25755_ (.A0(\cpuregs[10][14] ),
    .A1(_05121_),
    .S(_05603_),
    .X(_05606_));
 sky130_fd_sc_hd__clkbuf_1 _25756_ (.A(_05606_),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _25757_ (.A0(\cpuregs[10][15] ),
    .A1(_05129_),
    .S(_05603_),
    .X(_05607_));
 sky130_fd_sc_hd__clkbuf_1 _25758_ (.A(_05607_),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _25759_ (.A0(\cpuregs[10][16] ),
    .A1(_05138_),
    .S(_05603_),
    .X(_05608_));
 sky130_fd_sc_hd__clkbuf_1 _25760_ (.A(_05608_),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _25761_ (.A0(\cpuregs[10][17] ),
    .A1(_05146_),
    .S(_05603_),
    .X(_05609_));
 sky130_fd_sc_hd__clkbuf_1 _25762_ (.A(_05609_),
    .X(_00373_));
 sky130_fd_sc_hd__buf_2 _25763_ (.A(_05588_),
    .X(_05610_));
 sky130_fd_sc_hd__mux2_1 _25764_ (.A0(\cpuregs[10][18] ),
    .A1(_05154_),
    .S(_05610_),
    .X(_05611_));
 sky130_fd_sc_hd__clkbuf_1 _25765_ (.A(_05611_),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_1 _25766_ (.A0(\cpuregs[10][19] ),
    .A1(_05165_),
    .S(_05610_),
    .X(_05612_));
 sky130_fd_sc_hd__clkbuf_1 _25767_ (.A(_05612_),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _25768_ (.A0(\cpuregs[10][20] ),
    .A1(_05173_),
    .S(_05610_),
    .X(_05613_));
 sky130_fd_sc_hd__clkbuf_1 _25769_ (.A(_05613_),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _25770_ (.A0(\cpuregs[10][21] ),
    .A1(_05182_),
    .S(_05610_),
    .X(_05614_));
 sky130_fd_sc_hd__clkbuf_1 _25771_ (.A(_05614_),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_1 _25772_ (.A0(\cpuregs[10][22] ),
    .A1(_05191_),
    .S(_05610_),
    .X(_05615_));
 sky130_fd_sc_hd__clkbuf_1 _25773_ (.A(_05615_),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _25774_ (.A0(\cpuregs[10][23] ),
    .A1(_05199_),
    .S(_05610_),
    .X(_05616_));
 sky130_fd_sc_hd__clkbuf_1 _25775_ (.A(_05616_),
    .X(_00379_));
 sky130_fd_sc_hd__buf_2 _25776_ (.A(_05587_),
    .X(_05617_));
 sky130_fd_sc_hd__mux2_1 _25777_ (.A0(\cpuregs[10][24] ),
    .A1(_05206_),
    .S(_05617_),
    .X(_05618_));
 sky130_fd_sc_hd__clkbuf_1 _25778_ (.A(_05618_),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _25779_ (.A0(\cpuregs[10][25] ),
    .A1(_05217_),
    .S(_05617_),
    .X(_05619_));
 sky130_fd_sc_hd__clkbuf_1 _25780_ (.A(_05619_),
    .X(_00381_));
 sky130_fd_sc_hd__mux2_1 _25781_ (.A0(\cpuregs[10][26] ),
    .A1(_05225_),
    .S(_05617_),
    .X(_05620_));
 sky130_fd_sc_hd__clkbuf_1 _25782_ (.A(_05620_),
    .X(_00382_));
 sky130_fd_sc_hd__mux2_1 _25783_ (.A0(\cpuregs[10][27] ),
    .A1(_05232_),
    .S(_05617_),
    .X(_05621_));
 sky130_fd_sc_hd__clkbuf_1 _25784_ (.A(_05621_),
    .X(_00383_));
 sky130_fd_sc_hd__mux2_1 _25785_ (.A0(\cpuregs[10][28] ),
    .A1(_05240_),
    .S(_05617_),
    .X(_05622_));
 sky130_fd_sc_hd__clkbuf_1 _25786_ (.A(_05622_),
    .X(_00384_));
 sky130_fd_sc_hd__mux2_1 _25787_ (.A0(\cpuregs[10][29] ),
    .A1(_05248_),
    .S(_05617_),
    .X(_05623_));
 sky130_fd_sc_hd__clkbuf_1 _25788_ (.A(_05623_),
    .X(_00385_));
 sky130_fd_sc_hd__mux2_1 _25789_ (.A0(\cpuregs[10][30] ),
    .A1(_05256_),
    .S(_05588_),
    .X(_05624_));
 sky130_fd_sc_hd__clkbuf_1 _25790_ (.A(_05624_),
    .X(_00386_));
 sky130_fd_sc_hd__mux2_1 _25791_ (.A0(\cpuregs[10][31] ),
    .A1(_05263_),
    .S(_05588_),
    .X(_05625_));
 sky130_fd_sc_hd__clkbuf_1 _25792_ (.A(_05625_),
    .X(_00387_));
 sky130_fd_sc_hd__or2_1 _25793_ (.A(_05268_),
    .B(_05468_),
    .X(_05626_));
 sky130_fd_sc_hd__buf_4 _25794_ (.A(_05626_),
    .X(_05627_));
 sky130_fd_sc_hd__clkbuf_4 _25795_ (.A(_05627_),
    .X(_05628_));
 sky130_fd_sc_hd__mux2_1 _25796_ (.A0(_05265_),
    .A1(\cpuregs[11][0] ),
    .S(_05628_),
    .X(_05629_));
 sky130_fd_sc_hd__clkbuf_1 _25797_ (.A(_05629_),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _25798_ (.A0(_05274_),
    .A1(\cpuregs[11][1] ),
    .S(_05628_),
    .X(_05630_));
 sky130_fd_sc_hd__clkbuf_1 _25799_ (.A(_05630_),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_1 _25800_ (.A0(_05276_),
    .A1(\cpuregs[11][2] ),
    .S(_05628_),
    .X(_05631_));
 sky130_fd_sc_hd__clkbuf_1 _25801_ (.A(_05631_),
    .X(_00390_));
 sky130_fd_sc_hd__mux2_1 _25802_ (.A0(_05278_),
    .A1(\cpuregs[11][3] ),
    .S(_05628_),
    .X(_05632_));
 sky130_fd_sc_hd__clkbuf_1 _25803_ (.A(_05632_),
    .X(_00391_));
 sky130_fd_sc_hd__mux2_1 _25804_ (.A0(_05280_),
    .A1(\cpuregs[11][4] ),
    .S(_05628_),
    .X(_05633_));
 sky130_fd_sc_hd__clkbuf_1 _25805_ (.A(_05633_),
    .X(_00392_));
 sky130_fd_sc_hd__mux2_1 _25806_ (.A0(_05282_),
    .A1(\cpuregs[11][5] ),
    .S(_05628_),
    .X(_05634_));
 sky130_fd_sc_hd__clkbuf_1 _25807_ (.A(_05634_),
    .X(_00393_));
 sky130_fd_sc_hd__buf_2 _25808_ (.A(_05627_),
    .X(_05635_));
 sky130_fd_sc_hd__mux2_1 _25809_ (.A0(_05284_),
    .A1(\cpuregs[11][6] ),
    .S(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__clkbuf_1 _25810_ (.A(_05636_),
    .X(_00394_));
 sky130_fd_sc_hd__mux2_1 _25811_ (.A0(_05287_),
    .A1(\cpuregs[11][7] ),
    .S(_05635_),
    .X(_05637_));
 sky130_fd_sc_hd__clkbuf_1 _25812_ (.A(_05637_),
    .X(_00395_));
 sky130_fd_sc_hd__mux2_1 _25813_ (.A0(_05289_),
    .A1(\cpuregs[11][8] ),
    .S(_05635_),
    .X(_05638_));
 sky130_fd_sc_hd__clkbuf_1 _25814_ (.A(_05638_),
    .X(_00396_));
 sky130_fd_sc_hd__mux2_1 _25815_ (.A0(_05291_),
    .A1(\cpuregs[11][9] ),
    .S(_05635_),
    .X(_05639_));
 sky130_fd_sc_hd__clkbuf_1 _25816_ (.A(_05639_),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_1 _25817_ (.A0(_05293_),
    .A1(\cpuregs[11][10] ),
    .S(_05635_),
    .X(_05640_));
 sky130_fd_sc_hd__clkbuf_1 _25818_ (.A(_05640_),
    .X(_00398_));
 sky130_fd_sc_hd__mux2_1 _25819_ (.A0(_05295_),
    .A1(\cpuregs[11][11] ),
    .S(_05635_),
    .X(_05641_));
 sky130_fd_sc_hd__clkbuf_1 _25820_ (.A(_05641_),
    .X(_00399_));
 sky130_fd_sc_hd__buf_2 _25821_ (.A(_05627_),
    .X(_05642_));
 sky130_fd_sc_hd__mux2_1 _25822_ (.A0(_05297_),
    .A1(\cpuregs[11][12] ),
    .S(_05642_),
    .X(_05643_));
 sky130_fd_sc_hd__clkbuf_1 _25823_ (.A(_05643_),
    .X(_00400_));
 sky130_fd_sc_hd__mux2_1 _25824_ (.A0(_05300_),
    .A1(\cpuregs[11][13] ),
    .S(_05642_),
    .X(_05644_));
 sky130_fd_sc_hd__clkbuf_1 _25825_ (.A(_05644_),
    .X(_00401_));
 sky130_fd_sc_hd__mux2_1 _25826_ (.A0(_05302_),
    .A1(\cpuregs[11][14] ),
    .S(_05642_),
    .X(_05645_));
 sky130_fd_sc_hd__clkbuf_1 _25827_ (.A(_05645_),
    .X(_00402_));
 sky130_fd_sc_hd__mux2_1 _25828_ (.A0(_05304_),
    .A1(\cpuregs[11][15] ),
    .S(_05642_),
    .X(_05646_));
 sky130_fd_sc_hd__clkbuf_1 _25829_ (.A(_05646_),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _25830_ (.A0(_05306_),
    .A1(\cpuregs[11][16] ),
    .S(_05642_),
    .X(_05647_));
 sky130_fd_sc_hd__clkbuf_1 _25831_ (.A(_05647_),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_1 _25832_ (.A0(_05308_),
    .A1(\cpuregs[11][17] ),
    .S(_05642_),
    .X(_05648_));
 sky130_fd_sc_hd__clkbuf_1 _25833_ (.A(_05648_),
    .X(_00405_));
 sky130_fd_sc_hd__clkbuf_2 _25834_ (.A(_05627_),
    .X(_05649_));
 sky130_fd_sc_hd__mux2_1 _25835_ (.A0(_05310_),
    .A1(\cpuregs[11][18] ),
    .S(_05649_),
    .X(_05650_));
 sky130_fd_sc_hd__clkbuf_1 _25836_ (.A(_05650_),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_1 _25837_ (.A0(_05313_),
    .A1(\cpuregs[11][19] ),
    .S(_05649_),
    .X(_05651_));
 sky130_fd_sc_hd__clkbuf_1 _25838_ (.A(_05651_),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_1 _25839_ (.A0(_05315_),
    .A1(\cpuregs[11][20] ),
    .S(_05649_),
    .X(_05652_));
 sky130_fd_sc_hd__clkbuf_1 _25840_ (.A(_05652_),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_1 _25841_ (.A0(_05317_),
    .A1(\cpuregs[11][21] ),
    .S(_05649_),
    .X(_05653_));
 sky130_fd_sc_hd__clkbuf_1 _25842_ (.A(_05653_),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_1 _25843_ (.A0(_05319_),
    .A1(\cpuregs[11][22] ),
    .S(_05649_),
    .X(_05654_));
 sky130_fd_sc_hd__clkbuf_1 _25844_ (.A(_05654_),
    .X(_00410_));
 sky130_fd_sc_hd__mux2_1 _25845_ (.A0(_05321_),
    .A1(\cpuregs[11][23] ),
    .S(_05649_),
    .X(_05655_));
 sky130_fd_sc_hd__clkbuf_1 _25846_ (.A(_05655_),
    .X(_00411_));
 sky130_fd_sc_hd__clkbuf_4 _25847_ (.A(_05626_),
    .X(_05656_));
 sky130_fd_sc_hd__mux2_1 _25848_ (.A0(_05323_),
    .A1(\cpuregs[11][24] ),
    .S(_05656_),
    .X(_05657_));
 sky130_fd_sc_hd__clkbuf_1 _25849_ (.A(_05657_),
    .X(_00412_));
 sky130_fd_sc_hd__mux2_1 _25850_ (.A0(_05326_),
    .A1(\cpuregs[11][25] ),
    .S(_05656_),
    .X(_05658_));
 sky130_fd_sc_hd__clkbuf_1 _25851_ (.A(_05658_),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _25852_ (.A0(_05328_),
    .A1(\cpuregs[11][26] ),
    .S(_05656_),
    .X(_05659_));
 sky130_fd_sc_hd__clkbuf_1 _25853_ (.A(_05659_),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_1 _25854_ (.A0(_05330_),
    .A1(\cpuregs[11][27] ),
    .S(_05656_),
    .X(_05660_));
 sky130_fd_sc_hd__clkbuf_1 _25855_ (.A(_05660_),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _25856_ (.A0(_05332_),
    .A1(\cpuregs[11][28] ),
    .S(_05656_),
    .X(_05661_));
 sky130_fd_sc_hd__clkbuf_1 _25857_ (.A(_05661_),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _25858_ (.A0(_05334_),
    .A1(\cpuregs[11][29] ),
    .S(_05656_),
    .X(_05662_));
 sky130_fd_sc_hd__clkbuf_1 _25859_ (.A(_05662_),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _25860_ (.A0(_05336_),
    .A1(\cpuregs[11][30] ),
    .S(_05627_),
    .X(_05663_));
 sky130_fd_sc_hd__clkbuf_1 _25861_ (.A(_05663_),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _25862_ (.A0(_05338_),
    .A1(\cpuregs[11][31] ),
    .S(_05627_),
    .X(_05664_));
 sky130_fd_sc_hd__clkbuf_1 _25863_ (.A(_05664_),
    .X(_00419_));
 sky130_fd_sc_hd__clkbuf_2 _25864_ (.A(_04987_),
    .X(_05665_));
 sky130_fd_sc_hd__nand3b_1 _25865_ (.A_N(\latched_rd[4] ),
    .B(\latched_rd[3] ),
    .C(\latched_rd[2] ),
    .Y(_05666_));
 sky130_fd_sc_hd__nor2_1 _25866_ (.A(_04990_),
    .B(_05666_),
    .Y(_05667_));
 sky130_fd_sc_hd__buf_4 _25867_ (.A(_05667_),
    .X(_05668_));
 sky130_fd_sc_hd__buf_2 _25868_ (.A(_05668_),
    .X(_05669_));
 sky130_fd_sc_hd__mux2_1 _25869_ (.A0(\cpuregs[12][0] ),
    .A1(_05665_),
    .S(_05669_),
    .X(_05670_));
 sky130_fd_sc_hd__clkbuf_1 _25870_ (.A(_05670_),
    .X(_00420_));
 sky130_fd_sc_hd__clkbuf_2 _25871_ (.A(_05005_),
    .X(_05671_));
 sky130_fd_sc_hd__mux2_1 _25872_ (.A0(\cpuregs[12][1] ),
    .A1(_05671_),
    .S(_05669_),
    .X(_05672_));
 sky130_fd_sc_hd__clkbuf_1 _25873_ (.A(_05672_),
    .X(_00421_));
 sky130_fd_sc_hd__clkbuf_2 _25874_ (.A(_05015_),
    .X(_05673_));
 sky130_fd_sc_hd__mux2_1 _25875_ (.A0(\cpuregs[12][2] ),
    .A1(_05673_),
    .S(_05669_),
    .X(_05674_));
 sky130_fd_sc_hd__clkbuf_1 _25876_ (.A(_05674_),
    .X(_00422_));
 sky130_fd_sc_hd__buf_2 _25877_ (.A(_05022_),
    .X(_05675_));
 sky130_fd_sc_hd__mux2_1 _25878_ (.A0(\cpuregs[12][3] ),
    .A1(_05675_),
    .S(_05669_),
    .X(_05676_));
 sky130_fd_sc_hd__clkbuf_1 _25879_ (.A(_05676_),
    .X(_00423_));
 sky130_fd_sc_hd__buf_2 _25880_ (.A(_05031_),
    .X(_05677_));
 sky130_fd_sc_hd__mux2_1 _25881_ (.A0(\cpuregs[12][4] ),
    .A1(_05677_),
    .S(_05669_),
    .X(_05678_));
 sky130_fd_sc_hd__clkbuf_1 _25882_ (.A(_05678_),
    .X(_00424_));
 sky130_fd_sc_hd__clkbuf_2 _25883_ (.A(_05040_),
    .X(_05679_));
 sky130_fd_sc_hd__mux2_1 _25884_ (.A0(\cpuregs[12][5] ),
    .A1(_05679_),
    .S(_05669_),
    .X(_05680_));
 sky130_fd_sc_hd__clkbuf_1 _25885_ (.A(_05680_),
    .X(_00425_));
 sky130_fd_sc_hd__buf_2 _25886_ (.A(_05048_),
    .X(_05681_));
 sky130_fd_sc_hd__clkbuf_4 _25887_ (.A(_05668_),
    .X(_05682_));
 sky130_fd_sc_hd__mux2_1 _25888_ (.A0(\cpuregs[12][6] ),
    .A1(_05681_),
    .S(_05682_),
    .X(_05683_));
 sky130_fd_sc_hd__clkbuf_1 _25889_ (.A(_05683_),
    .X(_00426_));
 sky130_fd_sc_hd__clkbuf_4 _25890_ (.A(_05059_),
    .X(_05684_));
 sky130_fd_sc_hd__mux2_1 _25891_ (.A0(\cpuregs[12][7] ),
    .A1(_05684_),
    .S(_05682_),
    .X(_05685_));
 sky130_fd_sc_hd__clkbuf_1 _25892_ (.A(_05685_),
    .X(_00427_));
 sky130_fd_sc_hd__clkbuf_4 _25893_ (.A(_05068_),
    .X(_05686_));
 sky130_fd_sc_hd__mux2_1 _25894_ (.A0(\cpuregs[12][8] ),
    .A1(_05686_),
    .S(_05682_),
    .X(_05687_));
 sky130_fd_sc_hd__clkbuf_1 _25895_ (.A(_05687_),
    .X(_00428_));
 sky130_fd_sc_hd__buf_2 _25896_ (.A(_05075_),
    .X(_05688_));
 sky130_fd_sc_hd__mux2_1 _25897_ (.A0(\cpuregs[12][9] ),
    .A1(_05688_),
    .S(_05682_),
    .X(_05689_));
 sky130_fd_sc_hd__clkbuf_1 _25898_ (.A(_05689_),
    .X(_00429_));
 sky130_fd_sc_hd__clkbuf_4 _25899_ (.A(_05084_),
    .X(_05690_));
 sky130_fd_sc_hd__mux2_1 _25900_ (.A0(\cpuregs[12][10] ),
    .A1(_05690_),
    .S(_05682_),
    .X(_05691_));
 sky130_fd_sc_hd__clkbuf_1 _25901_ (.A(_05691_),
    .X(_00430_));
 sky130_fd_sc_hd__buf_2 _25902_ (.A(_05094_),
    .X(_05692_));
 sky130_fd_sc_hd__mux2_1 _25903_ (.A0(\cpuregs[12][11] ),
    .A1(_05692_),
    .S(_05682_),
    .X(_05693_));
 sky130_fd_sc_hd__clkbuf_1 _25904_ (.A(_05693_),
    .X(_00431_));
 sky130_fd_sc_hd__buf_2 _25905_ (.A(_05101_),
    .X(_05694_));
 sky130_fd_sc_hd__buf_2 _25906_ (.A(_05668_),
    .X(_05695_));
 sky130_fd_sc_hd__mux2_1 _25907_ (.A0(\cpuregs[12][12] ),
    .A1(_05694_),
    .S(_05695_),
    .X(_05696_));
 sky130_fd_sc_hd__clkbuf_1 _25908_ (.A(_05696_),
    .X(_00432_));
 sky130_fd_sc_hd__clkbuf_2 _25909_ (.A(_05112_),
    .X(_05697_));
 sky130_fd_sc_hd__mux2_1 _25910_ (.A0(\cpuregs[12][13] ),
    .A1(_05697_),
    .S(_05695_),
    .X(_05698_));
 sky130_fd_sc_hd__clkbuf_1 _25911_ (.A(_05698_),
    .X(_00433_));
 sky130_fd_sc_hd__clkbuf_2 _25912_ (.A(_05120_),
    .X(_05699_));
 sky130_fd_sc_hd__mux2_1 _25913_ (.A0(\cpuregs[12][14] ),
    .A1(_05699_),
    .S(_05695_),
    .X(_05700_));
 sky130_fd_sc_hd__clkbuf_1 _25914_ (.A(_05700_),
    .X(_00434_));
 sky130_fd_sc_hd__buf_2 _25915_ (.A(_05128_),
    .X(_05701_));
 sky130_fd_sc_hd__mux2_1 _25916_ (.A0(\cpuregs[12][15] ),
    .A1(_05701_),
    .S(_05695_),
    .X(_05702_));
 sky130_fd_sc_hd__clkbuf_1 _25917_ (.A(_05702_),
    .X(_00435_));
 sky130_fd_sc_hd__buf_2 _25918_ (.A(_05137_),
    .X(_05703_));
 sky130_fd_sc_hd__mux2_1 _25919_ (.A0(\cpuregs[12][16] ),
    .A1(_05703_),
    .S(_05695_),
    .X(_05704_));
 sky130_fd_sc_hd__clkbuf_1 _25920_ (.A(_05704_),
    .X(_00436_));
 sky130_fd_sc_hd__clkbuf_2 _25921_ (.A(_05145_),
    .X(_05705_));
 sky130_fd_sc_hd__mux2_1 _25922_ (.A0(\cpuregs[12][17] ),
    .A1(_05705_),
    .S(_05695_),
    .X(_05706_));
 sky130_fd_sc_hd__clkbuf_1 _25923_ (.A(_05706_),
    .X(_00437_));
 sky130_fd_sc_hd__clkbuf_2 _25924_ (.A(_05153_),
    .X(_05707_));
 sky130_fd_sc_hd__buf_2 _25925_ (.A(_05668_),
    .X(_05708_));
 sky130_fd_sc_hd__mux2_1 _25926_ (.A0(\cpuregs[12][18] ),
    .A1(_05707_),
    .S(_05708_),
    .X(_05709_));
 sky130_fd_sc_hd__clkbuf_1 _25927_ (.A(_05709_),
    .X(_00438_));
 sky130_fd_sc_hd__buf_2 _25928_ (.A(_05164_),
    .X(_05710_));
 sky130_fd_sc_hd__mux2_1 _25929_ (.A0(\cpuregs[12][19] ),
    .A1(_05710_),
    .S(_05708_),
    .X(_05711_));
 sky130_fd_sc_hd__clkbuf_1 _25930_ (.A(_05711_),
    .X(_00439_));
 sky130_fd_sc_hd__clkbuf_2 _25931_ (.A(_05172_),
    .X(_05712_));
 sky130_fd_sc_hd__mux2_1 _25932_ (.A0(\cpuregs[12][20] ),
    .A1(_05712_),
    .S(_05708_),
    .X(_05713_));
 sky130_fd_sc_hd__clkbuf_1 _25933_ (.A(_05713_),
    .X(_00440_));
 sky130_fd_sc_hd__buf_2 _25934_ (.A(_05181_),
    .X(_05714_));
 sky130_fd_sc_hd__mux2_1 _25935_ (.A0(\cpuregs[12][21] ),
    .A1(_05714_),
    .S(_05708_),
    .X(_05715_));
 sky130_fd_sc_hd__clkbuf_1 _25936_ (.A(_05715_),
    .X(_00441_));
 sky130_fd_sc_hd__clkbuf_2 _25937_ (.A(_05190_),
    .X(_05716_));
 sky130_fd_sc_hd__mux2_1 _25938_ (.A0(\cpuregs[12][22] ),
    .A1(_05716_),
    .S(_05708_),
    .X(_05717_));
 sky130_fd_sc_hd__clkbuf_1 _25939_ (.A(_05717_),
    .X(_00442_));
 sky130_fd_sc_hd__clkbuf_2 _25940_ (.A(_05198_),
    .X(_05718_));
 sky130_fd_sc_hd__mux2_1 _25941_ (.A0(\cpuregs[12][23] ),
    .A1(_05718_),
    .S(_05708_),
    .X(_05719_));
 sky130_fd_sc_hd__clkbuf_1 _25942_ (.A(_05719_),
    .X(_00443_));
 sky130_fd_sc_hd__buf_2 _25943_ (.A(_05205_),
    .X(_05720_));
 sky130_fd_sc_hd__clkbuf_4 _25944_ (.A(_05667_),
    .X(_05721_));
 sky130_fd_sc_hd__mux2_1 _25945_ (.A0(\cpuregs[12][24] ),
    .A1(_05720_),
    .S(_05721_),
    .X(_05722_));
 sky130_fd_sc_hd__clkbuf_1 _25946_ (.A(_05722_),
    .X(_00444_));
 sky130_fd_sc_hd__buf_2 _25947_ (.A(_05216_),
    .X(_05723_));
 sky130_fd_sc_hd__mux2_1 _25948_ (.A0(\cpuregs[12][25] ),
    .A1(_05723_),
    .S(_05721_),
    .X(_05724_));
 sky130_fd_sc_hd__clkbuf_1 _25949_ (.A(_05724_),
    .X(_00445_));
 sky130_fd_sc_hd__buf_2 _25950_ (.A(_05224_),
    .X(_05725_));
 sky130_fd_sc_hd__mux2_1 _25951_ (.A0(\cpuregs[12][26] ),
    .A1(_05725_),
    .S(_05721_),
    .X(_05726_));
 sky130_fd_sc_hd__clkbuf_1 _25952_ (.A(_05726_),
    .X(_00446_));
 sky130_fd_sc_hd__clkbuf_2 _25953_ (.A(_05231_),
    .X(_05727_));
 sky130_fd_sc_hd__mux2_1 _25954_ (.A0(\cpuregs[12][27] ),
    .A1(_05727_),
    .S(_05721_),
    .X(_05728_));
 sky130_fd_sc_hd__clkbuf_1 _25955_ (.A(_05728_),
    .X(_00447_));
 sky130_fd_sc_hd__clkbuf_2 _25956_ (.A(_05239_),
    .X(_05729_));
 sky130_fd_sc_hd__mux2_1 _25957_ (.A0(\cpuregs[12][28] ),
    .A1(_05729_),
    .S(_05721_),
    .X(_05730_));
 sky130_fd_sc_hd__clkbuf_1 _25958_ (.A(_05730_),
    .X(_00448_));
 sky130_fd_sc_hd__clkbuf_2 _25959_ (.A(_05247_),
    .X(_05731_));
 sky130_fd_sc_hd__mux2_1 _25960_ (.A0(\cpuregs[12][29] ),
    .A1(_05731_),
    .S(_05721_),
    .X(_05732_));
 sky130_fd_sc_hd__clkbuf_1 _25961_ (.A(_05732_),
    .X(_00449_));
 sky130_fd_sc_hd__buf_2 _25962_ (.A(_05255_),
    .X(_05733_));
 sky130_fd_sc_hd__mux2_1 _25963_ (.A0(\cpuregs[12][30] ),
    .A1(_05733_),
    .S(_05668_),
    .X(_05734_));
 sky130_fd_sc_hd__clkbuf_1 _25964_ (.A(_05734_),
    .X(_00450_));
 sky130_fd_sc_hd__buf_2 _25965_ (.A(_05262_),
    .X(_05735_));
 sky130_fd_sc_hd__mux2_1 _25966_ (.A0(\cpuregs[12][31] ),
    .A1(_05735_),
    .S(_05668_),
    .X(_05736_));
 sky130_fd_sc_hd__clkbuf_1 _25967_ (.A(_05736_),
    .X(_00451_));
 sky130_fd_sc_hd__nor2_1 _25968_ (.A(_08170_),
    .B(net332),
    .Y(_05737_));
 sky130_fd_sc_hd__or2_2 _25969_ (.A(_08170_),
    .B(net332),
    .X(_05738_));
 sky130_fd_sc_hd__or3_1 _25970_ (.A(_08163_),
    .B(\mem_state[1] ),
    .C(\mem_state[0] ),
    .X(_05739_));
 sky130_fd_sc_hd__or3b_1 _25971_ (.A(_08156_),
    .B(_08154_),
    .C_N(_05509_),
    .X(_05740_));
 sky130_fd_sc_hd__o31a_1 _25972_ (.A1(_08151_),
    .A2(_10341_),
    .A3(_05739_),
    .B1(_05740_),
    .X(_05741_));
 sky130_fd_sc_hd__nand2_1 _25973_ (.A(_08328_),
    .B(net332),
    .Y(_05742_));
 sky130_fd_sc_hd__o22a_1 _25974_ (.A1(_05738_),
    .A2(_05741_),
    .B1(_05742_),
    .B2(net65),
    .X(_05743_));
 sky130_fd_sc_hd__a21bo_1 _25975_ (.A1(_08156_),
    .A2(_05737_),
    .B1_N(_05743_),
    .X(_05744_));
 sky130_fd_sc_hd__and3_2 _25976_ (.A(mem_do_wdata),
    .B(_08154_),
    .C(_05737_),
    .X(_05745_));
 sky130_fd_sc_hd__o21bai_4 _25977_ (.A1(_08524_),
    .A2(_05738_),
    .B1_N(_05745_),
    .Y(_05746_));
 sky130_fd_sc_hd__buf_2 _25978_ (.A(_05746_),
    .X(_05747_));
 sky130_fd_sc_hd__clkbuf_4 _25979_ (.A(_05747_),
    .X(_05748_));
 sky130_fd_sc_hd__a21o_1 _25980_ (.A1(net198),
    .A2(_05744_),
    .B1(_05748_),
    .X(_00452_));
 sky130_fd_sc_hd__or2_1 _25981_ (.A(_05340_),
    .B(_05666_),
    .X(_05749_));
 sky130_fd_sc_hd__clkbuf_4 _25982_ (.A(_05749_),
    .X(_05750_));
 sky130_fd_sc_hd__buf_2 _25983_ (.A(_05750_),
    .X(_05751_));
 sky130_fd_sc_hd__mux2_1 _25984_ (.A0(_05265_),
    .A1(\cpuregs[13][0] ),
    .S(_05751_),
    .X(_05752_));
 sky130_fd_sc_hd__clkbuf_1 _25985_ (.A(_05752_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _25986_ (.A0(_05274_),
    .A1(\cpuregs[13][1] ),
    .S(_05751_),
    .X(_05753_));
 sky130_fd_sc_hd__clkbuf_1 _25987_ (.A(_05753_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _25988_ (.A0(_05276_),
    .A1(\cpuregs[13][2] ),
    .S(_05751_),
    .X(_05754_));
 sky130_fd_sc_hd__clkbuf_1 _25989_ (.A(_05754_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _25990_ (.A0(_05278_),
    .A1(\cpuregs[13][3] ),
    .S(_05751_),
    .X(_05755_));
 sky130_fd_sc_hd__clkbuf_1 _25991_ (.A(_05755_),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _25992_ (.A0(_05280_),
    .A1(\cpuregs[13][4] ),
    .S(_05751_),
    .X(_05756_));
 sky130_fd_sc_hd__clkbuf_1 _25993_ (.A(_05756_),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _25994_ (.A0(_05282_),
    .A1(\cpuregs[13][5] ),
    .S(_05751_),
    .X(_05757_));
 sky130_fd_sc_hd__clkbuf_1 _25995_ (.A(_05757_),
    .X(_00458_));
 sky130_fd_sc_hd__clkbuf_4 _25996_ (.A(_05750_),
    .X(_05758_));
 sky130_fd_sc_hd__mux2_1 _25997_ (.A0(_05284_),
    .A1(\cpuregs[13][6] ),
    .S(_05758_),
    .X(_05759_));
 sky130_fd_sc_hd__clkbuf_1 _25998_ (.A(_05759_),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _25999_ (.A0(_05287_),
    .A1(\cpuregs[13][7] ),
    .S(_05758_),
    .X(_05760_));
 sky130_fd_sc_hd__clkbuf_1 _26000_ (.A(_05760_),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _26001_ (.A0(_05289_),
    .A1(\cpuregs[13][8] ),
    .S(_05758_),
    .X(_05761_));
 sky130_fd_sc_hd__clkbuf_1 _26002_ (.A(_05761_),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _26003_ (.A0(_05291_),
    .A1(\cpuregs[13][9] ),
    .S(_05758_),
    .X(_05762_));
 sky130_fd_sc_hd__clkbuf_1 _26004_ (.A(_05762_),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _26005_ (.A0(_05293_),
    .A1(\cpuregs[13][10] ),
    .S(_05758_),
    .X(_05763_));
 sky130_fd_sc_hd__clkbuf_1 _26006_ (.A(_05763_),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _26007_ (.A0(_05295_),
    .A1(\cpuregs[13][11] ),
    .S(_05758_),
    .X(_05764_));
 sky130_fd_sc_hd__clkbuf_1 _26008_ (.A(_05764_),
    .X(_00464_));
 sky130_fd_sc_hd__clkbuf_2 _26009_ (.A(_05750_),
    .X(_05765_));
 sky130_fd_sc_hd__mux2_1 _26010_ (.A0(_05297_),
    .A1(\cpuregs[13][12] ),
    .S(_05765_),
    .X(_05766_));
 sky130_fd_sc_hd__clkbuf_1 _26011_ (.A(_05766_),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _26012_ (.A0(_05300_),
    .A1(\cpuregs[13][13] ),
    .S(_05765_),
    .X(_05767_));
 sky130_fd_sc_hd__clkbuf_1 _26013_ (.A(_05767_),
    .X(_00466_));
 sky130_fd_sc_hd__mux2_1 _26014_ (.A0(_05302_),
    .A1(\cpuregs[13][14] ),
    .S(_05765_),
    .X(_05768_));
 sky130_fd_sc_hd__clkbuf_1 _26015_ (.A(_05768_),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _26016_ (.A0(_05304_),
    .A1(\cpuregs[13][15] ),
    .S(_05765_),
    .X(_05769_));
 sky130_fd_sc_hd__clkbuf_1 _26017_ (.A(_05769_),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _26018_ (.A0(_05306_),
    .A1(\cpuregs[13][16] ),
    .S(_05765_),
    .X(_05770_));
 sky130_fd_sc_hd__clkbuf_1 _26019_ (.A(_05770_),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _26020_ (.A0(_05308_),
    .A1(\cpuregs[13][17] ),
    .S(_05765_),
    .X(_05771_));
 sky130_fd_sc_hd__clkbuf_1 _26021_ (.A(_05771_),
    .X(_00470_));
 sky130_fd_sc_hd__buf_2 _26022_ (.A(_05750_),
    .X(_05772_));
 sky130_fd_sc_hd__mux2_1 _26023_ (.A0(_05310_),
    .A1(\cpuregs[13][18] ),
    .S(_05772_),
    .X(_05773_));
 sky130_fd_sc_hd__clkbuf_1 _26024_ (.A(_05773_),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _26025_ (.A0(_05313_),
    .A1(\cpuregs[13][19] ),
    .S(_05772_),
    .X(_05774_));
 sky130_fd_sc_hd__clkbuf_1 _26026_ (.A(_05774_),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _26027_ (.A0(_05315_),
    .A1(\cpuregs[13][20] ),
    .S(_05772_),
    .X(_05775_));
 sky130_fd_sc_hd__clkbuf_1 _26028_ (.A(_05775_),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _26029_ (.A0(_05317_),
    .A1(\cpuregs[13][21] ),
    .S(_05772_),
    .X(_05776_));
 sky130_fd_sc_hd__clkbuf_1 _26030_ (.A(_05776_),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _26031_ (.A0(_05319_),
    .A1(\cpuregs[13][22] ),
    .S(_05772_),
    .X(_05777_));
 sky130_fd_sc_hd__clkbuf_1 _26032_ (.A(_05777_),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _26033_ (.A0(_05321_),
    .A1(\cpuregs[13][23] ),
    .S(_05772_),
    .X(_05778_));
 sky130_fd_sc_hd__clkbuf_1 _26034_ (.A(_05778_),
    .X(_00476_));
 sky130_fd_sc_hd__clkbuf_4 _26035_ (.A(_05749_),
    .X(_05779_));
 sky130_fd_sc_hd__mux2_1 _26036_ (.A0(_05323_),
    .A1(\cpuregs[13][24] ),
    .S(_05779_),
    .X(_05780_));
 sky130_fd_sc_hd__clkbuf_1 _26037_ (.A(_05780_),
    .X(_00477_));
 sky130_fd_sc_hd__mux2_1 _26038_ (.A0(_05326_),
    .A1(\cpuregs[13][25] ),
    .S(_05779_),
    .X(_05781_));
 sky130_fd_sc_hd__clkbuf_1 _26039_ (.A(_05781_),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_1 _26040_ (.A0(_05328_),
    .A1(\cpuregs[13][26] ),
    .S(_05779_),
    .X(_05782_));
 sky130_fd_sc_hd__clkbuf_1 _26041_ (.A(_05782_),
    .X(_00479_));
 sky130_fd_sc_hd__mux2_1 _26042_ (.A0(_05330_),
    .A1(\cpuregs[13][27] ),
    .S(_05779_),
    .X(_05783_));
 sky130_fd_sc_hd__clkbuf_1 _26043_ (.A(_05783_),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_1 _26044_ (.A0(_05332_),
    .A1(\cpuregs[13][28] ),
    .S(_05779_),
    .X(_05784_));
 sky130_fd_sc_hd__clkbuf_1 _26045_ (.A(_05784_),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _26046_ (.A0(_05334_),
    .A1(\cpuregs[13][29] ),
    .S(_05779_),
    .X(_05785_));
 sky130_fd_sc_hd__clkbuf_1 _26047_ (.A(_05785_),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _26048_ (.A0(_05336_),
    .A1(\cpuregs[13][30] ),
    .S(_05750_),
    .X(_05786_));
 sky130_fd_sc_hd__clkbuf_1 _26049_ (.A(_05786_),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_1 _26050_ (.A0(_05338_),
    .A1(\cpuregs[13][31] ),
    .S(_05750_),
    .X(_05787_));
 sky130_fd_sc_hd__clkbuf_1 _26051_ (.A(_05787_),
    .X(_00484_));
 sky130_fd_sc_hd__or2_1 _26052_ (.A(_05381_),
    .B(_05666_),
    .X(_05788_));
 sky130_fd_sc_hd__buf_4 _26053_ (.A(_05788_),
    .X(_05789_));
 sky130_fd_sc_hd__buf_2 _26054_ (.A(_05789_),
    .X(_05790_));
 sky130_fd_sc_hd__mux2_1 _26055_ (.A0(_05265_),
    .A1(\cpuregs[14][0] ),
    .S(_05790_),
    .X(_05791_));
 sky130_fd_sc_hd__clkbuf_1 _26056_ (.A(_05791_),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _26057_ (.A0(_05274_),
    .A1(\cpuregs[14][1] ),
    .S(_05790_),
    .X(_05792_));
 sky130_fd_sc_hd__clkbuf_1 _26058_ (.A(_05792_),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _26059_ (.A0(_05276_),
    .A1(\cpuregs[14][2] ),
    .S(_05790_),
    .X(_05793_));
 sky130_fd_sc_hd__clkbuf_1 _26060_ (.A(_05793_),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _26061_ (.A0(_05278_),
    .A1(\cpuregs[14][3] ),
    .S(_05790_),
    .X(_05794_));
 sky130_fd_sc_hd__clkbuf_1 _26062_ (.A(_05794_),
    .X(_00488_));
 sky130_fd_sc_hd__mux2_1 _26063_ (.A0(_05280_),
    .A1(\cpuregs[14][4] ),
    .S(_05790_),
    .X(_05795_));
 sky130_fd_sc_hd__clkbuf_1 _26064_ (.A(_05795_),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_1 _26065_ (.A0(_05282_),
    .A1(\cpuregs[14][5] ),
    .S(_05790_),
    .X(_05796_));
 sky130_fd_sc_hd__clkbuf_1 _26066_ (.A(_05796_),
    .X(_00490_));
 sky130_fd_sc_hd__clkbuf_4 _26067_ (.A(_05789_),
    .X(_05797_));
 sky130_fd_sc_hd__mux2_1 _26068_ (.A0(_05284_),
    .A1(\cpuregs[14][6] ),
    .S(_05797_),
    .X(_05798_));
 sky130_fd_sc_hd__clkbuf_1 _26069_ (.A(_05798_),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_1 _26070_ (.A0(_05287_),
    .A1(\cpuregs[14][7] ),
    .S(_05797_),
    .X(_05799_));
 sky130_fd_sc_hd__clkbuf_1 _26071_ (.A(_05799_),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _26072_ (.A0(_05289_),
    .A1(\cpuregs[14][8] ),
    .S(_05797_),
    .X(_05800_));
 sky130_fd_sc_hd__clkbuf_1 _26073_ (.A(_05800_),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _26074_ (.A0(_05291_),
    .A1(\cpuregs[14][9] ),
    .S(_05797_),
    .X(_05801_));
 sky130_fd_sc_hd__clkbuf_1 _26075_ (.A(_05801_),
    .X(_00494_));
 sky130_fd_sc_hd__mux2_1 _26076_ (.A0(_05293_),
    .A1(\cpuregs[14][10] ),
    .S(_05797_),
    .X(_05802_));
 sky130_fd_sc_hd__clkbuf_1 _26077_ (.A(_05802_),
    .X(_00495_));
 sky130_fd_sc_hd__mux2_1 _26078_ (.A0(_05295_),
    .A1(\cpuregs[14][11] ),
    .S(_05797_),
    .X(_05803_));
 sky130_fd_sc_hd__clkbuf_1 _26079_ (.A(_05803_),
    .X(_00496_));
 sky130_fd_sc_hd__buf_2 _26080_ (.A(_05789_),
    .X(_05804_));
 sky130_fd_sc_hd__mux2_1 _26081_ (.A0(_05297_),
    .A1(\cpuregs[14][12] ),
    .S(_05804_),
    .X(_05805_));
 sky130_fd_sc_hd__clkbuf_1 _26082_ (.A(_05805_),
    .X(_00497_));
 sky130_fd_sc_hd__mux2_1 _26083_ (.A0(_05300_),
    .A1(\cpuregs[14][13] ),
    .S(_05804_),
    .X(_05806_));
 sky130_fd_sc_hd__clkbuf_1 _26084_ (.A(_05806_),
    .X(_00498_));
 sky130_fd_sc_hd__mux2_1 _26085_ (.A0(_05302_),
    .A1(\cpuregs[14][14] ),
    .S(_05804_),
    .X(_05807_));
 sky130_fd_sc_hd__clkbuf_1 _26086_ (.A(_05807_),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_1 _26087_ (.A0(_05304_),
    .A1(\cpuregs[14][15] ),
    .S(_05804_),
    .X(_05808_));
 sky130_fd_sc_hd__clkbuf_1 _26088_ (.A(_05808_),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _26089_ (.A0(_05306_),
    .A1(\cpuregs[14][16] ),
    .S(_05804_),
    .X(_05809_));
 sky130_fd_sc_hd__clkbuf_1 _26090_ (.A(_05809_),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _26091_ (.A0(_05308_),
    .A1(\cpuregs[14][17] ),
    .S(_05804_),
    .X(_05810_));
 sky130_fd_sc_hd__clkbuf_1 _26092_ (.A(_05810_),
    .X(_00502_));
 sky130_fd_sc_hd__clkbuf_2 _26093_ (.A(_05789_),
    .X(_05811_));
 sky130_fd_sc_hd__mux2_1 _26094_ (.A0(_05310_),
    .A1(\cpuregs[14][18] ),
    .S(_05811_),
    .X(_05812_));
 sky130_fd_sc_hd__clkbuf_1 _26095_ (.A(_05812_),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _26096_ (.A0(_05313_),
    .A1(\cpuregs[14][19] ),
    .S(_05811_),
    .X(_05813_));
 sky130_fd_sc_hd__clkbuf_1 _26097_ (.A(_05813_),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _26098_ (.A0(_05315_),
    .A1(\cpuregs[14][20] ),
    .S(_05811_),
    .X(_05814_));
 sky130_fd_sc_hd__clkbuf_1 _26099_ (.A(_05814_),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _26100_ (.A0(_05317_),
    .A1(\cpuregs[14][21] ),
    .S(_05811_),
    .X(_05815_));
 sky130_fd_sc_hd__clkbuf_1 _26101_ (.A(_05815_),
    .X(_00506_));
 sky130_fd_sc_hd__mux2_1 _26102_ (.A0(_05319_),
    .A1(\cpuregs[14][22] ),
    .S(_05811_),
    .X(_05816_));
 sky130_fd_sc_hd__clkbuf_1 _26103_ (.A(_05816_),
    .X(_00507_));
 sky130_fd_sc_hd__mux2_1 _26104_ (.A0(_05321_),
    .A1(\cpuregs[14][23] ),
    .S(_05811_),
    .X(_05817_));
 sky130_fd_sc_hd__clkbuf_1 _26105_ (.A(_05817_),
    .X(_00508_));
 sky130_fd_sc_hd__clkbuf_4 _26106_ (.A(_05788_),
    .X(_05818_));
 sky130_fd_sc_hd__mux2_1 _26107_ (.A0(_05323_),
    .A1(\cpuregs[14][24] ),
    .S(_05818_),
    .X(_05819_));
 sky130_fd_sc_hd__clkbuf_1 _26108_ (.A(_05819_),
    .X(_00509_));
 sky130_fd_sc_hd__mux2_1 _26109_ (.A0(_05326_),
    .A1(\cpuregs[14][25] ),
    .S(_05818_),
    .X(_05820_));
 sky130_fd_sc_hd__clkbuf_1 _26110_ (.A(_05820_),
    .X(_00510_));
 sky130_fd_sc_hd__mux2_1 _26111_ (.A0(_05328_),
    .A1(\cpuregs[14][26] ),
    .S(_05818_),
    .X(_05821_));
 sky130_fd_sc_hd__clkbuf_1 _26112_ (.A(_05821_),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _26113_ (.A0(_05330_),
    .A1(\cpuregs[14][27] ),
    .S(_05818_),
    .X(_05822_));
 sky130_fd_sc_hd__clkbuf_1 _26114_ (.A(_05822_),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_1 _26115_ (.A0(_05332_),
    .A1(\cpuregs[14][28] ),
    .S(_05818_),
    .X(_05823_));
 sky130_fd_sc_hd__clkbuf_1 _26116_ (.A(_05823_),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _26117_ (.A0(_05334_),
    .A1(\cpuregs[14][29] ),
    .S(_05818_),
    .X(_05824_));
 sky130_fd_sc_hd__clkbuf_1 _26118_ (.A(_05824_),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _26119_ (.A0(_05336_),
    .A1(\cpuregs[14][30] ),
    .S(_05789_),
    .X(_05825_));
 sky130_fd_sc_hd__clkbuf_1 _26120_ (.A(_05825_),
    .X(_00515_));
 sky130_fd_sc_hd__mux2_1 _26121_ (.A0(_05338_),
    .A1(\cpuregs[14][31] ),
    .S(_05789_),
    .X(_05826_));
 sky130_fd_sc_hd__clkbuf_1 _26122_ (.A(_05826_),
    .X(_00516_));
 sky130_fd_sc_hd__or2_1 _26123_ (.A(_05268_),
    .B(_05666_),
    .X(_05827_));
 sky130_fd_sc_hd__buf_4 _26124_ (.A(_05827_),
    .X(_05828_));
 sky130_fd_sc_hd__buf_2 _26125_ (.A(_05828_),
    .X(_05829_));
 sky130_fd_sc_hd__mux2_1 _26126_ (.A0(_05265_),
    .A1(\cpuregs[15][0] ),
    .S(_05829_),
    .X(_05830_));
 sky130_fd_sc_hd__clkbuf_1 _26127_ (.A(_05830_),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_1 _26128_ (.A0(_05274_),
    .A1(\cpuregs[15][1] ),
    .S(_05829_),
    .X(_05831_));
 sky130_fd_sc_hd__clkbuf_1 _26129_ (.A(_05831_),
    .X(_00518_));
 sky130_fd_sc_hd__mux2_1 _26130_ (.A0(_05276_),
    .A1(\cpuregs[15][2] ),
    .S(_05829_),
    .X(_05832_));
 sky130_fd_sc_hd__clkbuf_1 _26131_ (.A(_05832_),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_1 _26132_ (.A0(_05278_),
    .A1(\cpuregs[15][3] ),
    .S(_05829_),
    .X(_05833_));
 sky130_fd_sc_hd__clkbuf_1 _26133_ (.A(_05833_),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_1 _26134_ (.A0(_05280_),
    .A1(\cpuregs[15][4] ),
    .S(_05829_),
    .X(_05834_));
 sky130_fd_sc_hd__clkbuf_1 _26135_ (.A(_05834_),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _26136_ (.A0(_05282_),
    .A1(\cpuregs[15][5] ),
    .S(_05829_),
    .X(_05835_));
 sky130_fd_sc_hd__clkbuf_1 _26137_ (.A(_05835_),
    .X(_00522_));
 sky130_fd_sc_hd__buf_2 _26138_ (.A(_05828_),
    .X(_05836_));
 sky130_fd_sc_hd__mux2_1 _26139_ (.A0(_05284_),
    .A1(\cpuregs[15][6] ),
    .S(_05836_),
    .X(_05837_));
 sky130_fd_sc_hd__clkbuf_1 _26140_ (.A(_05837_),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _26141_ (.A0(_05287_),
    .A1(\cpuregs[15][7] ),
    .S(_05836_),
    .X(_05838_));
 sky130_fd_sc_hd__clkbuf_1 _26142_ (.A(_05838_),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _26143_ (.A0(_05289_),
    .A1(\cpuregs[15][8] ),
    .S(_05836_),
    .X(_05839_));
 sky130_fd_sc_hd__clkbuf_1 _26144_ (.A(_05839_),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_1 _26145_ (.A0(_05291_),
    .A1(\cpuregs[15][9] ),
    .S(_05836_),
    .X(_05840_));
 sky130_fd_sc_hd__clkbuf_1 _26146_ (.A(_05840_),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _26147_ (.A0(_05293_),
    .A1(\cpuregs[15][10] ),
    .S(_05836_),
    .X(_05841_));
 sky130_fd_sc_hd__clkbuf_1 _26148_ (.A(_05841_),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _26149_ (.A0(_05295_),
    .A1(\cpuregs[15][11] ),
    .S(_05836_),
    .X(_05842_));
 sky130_fd_sc_hd__clkbuf_1 _26150_ (.A(_05842_),
    .X(_00528_));
 sky130_fd_sc_hd__clkbuf_2 _26151_ (.A(_05828_),
    .X(_05843_));
 sky130_fd_sc_hd__mux2_1 _26152_ (.A0(_05297_),
    .A1(\cpuregs[15][12] ),
    .S(_05843_),
    .X(_05844_));
 sky130_fd_sc_hd__clkbuf_1 _26153_ (.A(_05844_),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_1 _26154_ (.A0(_05300_),
    .A1(\cpuregs[15][13] ),
    .S(_05843_),
    .X(_05845_));
 sky130_fd_sc_hd__clkbuf_1 _26155_ (.A(_05845_),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_1 _26156_ (.A0(_05302_),
    .A1(\cpuregs[15][14] ),
    .S(_05843_),
    .X(_05846_));
 sky130_fd_sc_hd__clkbuf_1 _26157_ (.A(_05846_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _26158_ (.A0(_05304_),
    .A1(\cpuregs[15][15] ),
    .S(_05843_),
    .X(_05847_));
 sky130_fd_sc_hd__clkbuf_1 _26159_ (.A(_05847_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _26160_ (.A0(_05306_),
    .A1(\cpuregs[15][16] ),
    .S(_05843_),
    .X(_05848_));
 sky130_fd_sc_hd__clkbuf_1 _26161_ (.A(_05848_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _26162_ (.A0(_05308_),
    .A1(\cpuregs[15][17] ),
    .S(_05843_),
    .X(_05849_));
 sky130_fd_sc_hd__clkbuf_1 _26163_ (.A(_05849_),
    .X(_00534_));
 sky130_fd_sc_hd__buf_2 _26164_ (.A(_05828_),
    .X(_05850_));
 sky130_fd_sc_hd__mux2_1 _26165_ (.A0(_05310_),
    .A1(\cpuregs[15][18] ),
    .S(_05850_),
    .X(_05851_));
 sky130_fd_sc_hd__clkbuf_1 _26166_ (.A(_05851_),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _26167_ (.A0(_05313_),
    .A1(\cpuregs[15][19] ),
    .S(_05850_),
    .X(_05852_));
 sky130_fd_sc_hd__clkbuf_1 _26168_ (.A(_05852_),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_1 _26169_ (.A0(_05315_),
    .A1(\cpuregs[15][20] ),
    .S(_05850_),
    .X(_05853_));
 sky130_fd_sc_hd__clkbuf_1 _26170_ (.A(_05853_),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_1 _26171_ (.A0(_05317_),
    .A1(\cpuregs[15][21] ),
    .S(_05850_),
    .X(_05854_));
 sky130_fd_sc_hd__clkbuf_1 _26172_ (.A(_05854_),
    .X(_00538_));
 sky130_fd_sc_hd__mux2_1 _26173_ (.A0(_05319_),
    .A1(\cpuregs[15][22] ),
    .S(_05850_),
    .X(_05855_));
 sky130_fd_sc_hd__clkbuf_1 _26174_ (.A(_05855_),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _26175_ (.A0(_05321_),
    .A1(\cpuregs[15][23] ),
    .S(_05850_),
    .X(_05856_));
 sky130_fd_sc_hd__clkbuf_1 _26176_ (.A(_05856_),
    .X(_00540_));
 sky130_fd_sc_hd__buf_2 _26177_ (.A(_05827_),
    .X(_05857_));
 sky130_fd_sc_hd__mux2_1 _26178_ (.A0(_05323_),
    .A1(\cpuregs[15][24] ),
    .S(_05857_),
    .X(_05858_));
 sky130_fd_sc_hd__clkbuf_1 _26179_ (.A(_05858_),
    .X(_00541_));
 sky130_fd_sc_hd__mux2_1 _26180_ (.A0(_05326_),
    .A1(\cpuregs[15][25] ),
    .S(_05857_),
    .X(_05859_));
 sky130_fd_sc_hd__clkbuf_1 _26181_ (.A(_05859_),
    .X(_00542_));
 sky130_fd_sc_hd__mux2_1 _26182_ (.A0(_05328_),
    .A1(\cpuregs[15][26] ),
    .S(_05857_),
    .X(_05860_));
 sky130_fd_sc_hd__clkbuf_1 _26183_ (.A(_05860_),
    .X(_00543_));
 sky130_fd_sc_hd__mux2_1 _26184_ (.A0(_05330_),
    .A1(\cpuregs[15][27] ),
    .S(_05857_),
    .X(_05861_));
 sky130_fd_sc_hd__clkbuf_1 _26185_ (.A(_05861_),
    .X(_00544_));
 sky130_fd_sc_hd__mux2_1 _26186_ (.A0(_05332_),
    .A1(\cpuregs[15][28] ),
    .S(_05857_),
    .X(_05862_));
 sky130_fd_sc_hd__clkbuf_1 _26187_ (.A(_05862_),
    .X(_00545_));
 sky130_fd_sc_hd__mux2_1 _26188_ (.A0(_05334_),
    .A1(\cpuregs[15][29] ),
    .S(_05857_),
    .X(_05863_));
 sky130_fd_sc_hd__clkbuf_1 _26189_ (.A(_05863_),
    .X(_00546_));
 sky130_fd_sc_hd__mux2_1 _26190_ (.A0(_05336_),
    .A1(\cpuregs[15][30] ),
    .S(_05828_),
    .X(_05864_));
 sky130_fd_sc_hd__clkbuf_1 _26191_ (.A(_05864_),
    .X(_00547_));
 sky130_fd_sc_hd__mux2_1 _26192_ (.A0(_05338_),
    .A1(\cpuregs[15][31] ),
    .S(_05828_),
    .X(_05865_));
 sky130_fd_sc_hd__clkbuf_1 _26193_ (.A(_05865_),
    .X(_00548_));
 sky130_fd_sc_hd__or3b_1 _26194_ (.A(\latched_rd[2] ),
    .B(\latched_rd[3] ),
    .C_N(\latched_rd[4] ),
    .X(_05866_));
 sky130_fd_sc_hd__nor2_1 _26195_ (.A(_04990_),
    .B(_05866_),
    .Y(_05867_));
 sky130_fd_sc_hd__clkbuf_2 _26196_ (.A(_05867_),
    .X(_05868_));
 sky130_fd_sc_hd__buf_2 _26197_ (.A(_05868_),
    .X(_05869_));
 sky130_fd_sc_hd__mux2_1 _26198_ (.A0(\cpuregs[16][0] ),
    .A1(_05665_),
    .S(_05869_),
    .X(_05870_));
 sky130_fd_sc_hd__clkbuf_1 _26199_ (.A(_05870_),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _26200_ (.A0(\cpuregs[16][1] ),
    .A1(_05671_),
    .S(_05869_),
    .X(_05871_));
 sky130_fd_sc_hd__clkbuf_1 _26201_ (.A(_05871_),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _26202_ (.A0(\cpuregs[16][2] ),
    .A1(_05673_),
    .S(_05869_),
    .X(_05872_));
 sky130_fd_sc_hd__clkbuf_1 _26203_ (.A(_05872_),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _26204_ (.A0(\cpuregs[16][3] ),
    .A1(_05675_),
    .S(_05869_),
    .X(_05873_));
 sky130_fd_sc_hd__clkbuf_1 _26205_ (.A(_05873_),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _26206_ (.A0(\cpuregs[16][4] ),
    .A1(_05677_),
    .S(_05869_),
    .X(_05874_));
 sky130_fd_sc_hd__clkbuf_1 _26207_ (.A(_05874_),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_1 _26208_ (.A0(\cpuregs[16][5] ),
    .A1(_05679_),
    .S(_05869_),
    .X(_05875_));
 sky130_fd_sc_hd__clkbuf_1 _26209_ (.A(_05875_),
    .X(_00554_));
 sky130_fd_sc_hd__buf_2 _26210_ (.A(_05868_),
    .X(_05876_));
 sky130_fd_sc_hd__mux2_1 _26211_ (.A0(\cpuregs[16][6] ),
    .A1(_05681_),
    .S(_05876_),
    .X(_05877_));
 sky130_fd_sc_hd__clkbuf_1 _26212_ (.A(_05877_),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_1 _26213_ (.A0(\cpuregs[16][7] ),
    .A1(_05684_),
    .S(_05876_),
    .X(_05878_));
 sky130_fd_sc_hd__clkbuf_1 _26214_ (.A(_05878_),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_1 _26215_ (.A0(\cpuregs[16][8] ),
    .A1(_05686_),
    .S(_05876_),
    .X(_05879_));
 sky130_fd_sc_hd__clkbuf_1 _26216_ (.A(_05879_),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _26217_ (.A0(\cpuregs[16][9] ),
    .A1(_05688_),
    .S(_05876_),
    .X(_05880_));
 sky130_fd_sc_hd__clkbuf_1 _26218_ (.A(_05880_),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_1 _26219_ (.A0(\cpuregs[16][10] ),
    .A1(_05690_),
    .S(_05876_),
    .X(_05881_));
 sky130_fd_sc_hd__clkbuf_1 _26220_ (.A(_05881_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _26221_ (.A0(\cpuregs[16][11] ),
    .A1(_05692_),
    .S(_05876_),
    .X(_05882_));
 sky130_fd_sc_hd__clkbuf_1 _26222_ (.A(_05882_),
    .X(_00560_));
 sky130_fd_sc_hd__buf_2 _26223_ (.A(_05868_),
    .X(_05883_));
 sky130_fd_sc_hd__mux2_1 _26224_ (.A0(\cpuregs[16][12] ),
    .A1(_05694_),
    .S(_05883_),
    .X(_05884_));
 sky130_fd_sc_hd__clkbuf_1 _26225_ (.A(_05884_),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _26226_ (.A0(\cpuregs[16][13] ),
    .A1(_05697_),
    .S(_05883_),
    .X(_05885_));
 sky130_fd_sc_hd__clkbuf_1 _26227_ (.A(_05885_),
    .X(_00562_));
 sky130_fd_sc_hd__mux2_1 _26228_ (.A0(\cpuregs[16][14] ),
    .A1(_05699_),
    .S(_05883_),
    .X(_05886_));
 sky130_fd_sc_hd__clkbuf_1 _26229_ (.A(_05886_),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _26230_ (.A0(\cpuregs[16][15] ),
    .A1(_05701_),
    .S(_05883_),
    .X(_05887_));
 sky130_fd_sc_hd__clkbuf_1 _26231_ (.A(_05887_),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _26232_ (.A0(\cpuregs[16][16] ),
    .A1(_05703_),
    .S(_05883_),
    .X(_05888_));
 sky130_fd_sc_hd__clkbuf_1 _26233_ (.A(_05888_),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _26234_ (.A0(\cpuregs[16][17] ),
    .A1(_05705_),
    .S(_05883_),
    .X(_05889_));
 sky130_fd_sc_hd__clkbuf_1 _26235_ (.A(_05889_),
    .X(_00566_));
 sky130_fd_sc_hd__buf_2 _26236_ (.A(_05868_),
    .X(_05890_));
 sky130_fd_sc_hd__mux2_1 _26237_ (.A0(\cpuregs[16][18] ),
    .A1(_05707_),
    .S(_05890_),
    .X(_05891_));
 sky130_fd_sc_hd__clkbuf_1 _26238_ (.A(_05891_),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _26239_ (.A0(\cpuregs[16][19] ),
    .A1(_05710_),
    .S(_05890_),
    .X(_05892_));
 sky130_fd_sc_hd__clkbuf_1 _26240_ (.A(_05892_),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _26241_ (.A0(\cpuregs[16][20] ),
    .A1(_05712_),
    .S(_05890_),
    .X(_05893_));
 sky130_fd_sc_hd__clkbuf_1 _26242_ (.A(_05893_),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _26243_ (.A0(\cpuregs[16][21] ),
    .A1(_05714_),
    .S(_05890_),
    .X(_05894_));
 sky130_fd_sc_hd__clkbuf_1 _26244_ (.A(_05894_),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _26245_ (.A0(\cpuregs[16][22] ),
    .A1(_05716_),
    .S(_05890_),
    .X(_05895_));
 sky130_fd_sc_hd__clkbuf_1 _26246_ (.A(_05895_),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_1 _26247_ (.A0(\cpuregs[16][23] ),
    .A1(_05718_),
    .S(_05890_),
    .X(_05896_));
 sky130_fd_sc_hd__clkbuf_1 _26248_ (.A(_05896_),
    .X(_00572_));
 sky130_fd_sc_hd__buf_2 _26249_ (.A(_05867_),
    .X(_05897_));
 sky130_fd_sc_hd__mux2_1 _26250_ (.A0(\cpuregs[16][24] ),
    .A1(_05720_),
    .S(_05897_),
    .X(_05898_));
 sky130_fd_sc_hd__clkbuf_1 _26251_ (.A(_05898_),
    .X(_00573_));
 sky130_fd_sc_hd__mux2_1 _26252_ (.A0(\cpuregs[16][25] ),
    .A1(_05723_),
    .S(_05897_),
    .X(_05899_));
 sky130_fd_sc_hd__clkbuf_1 _26253_ (.A(_05899_),
    .X(_00574_));
 sky130_fd_sc_hd__mux2_1 _26254_ (.A0(\cpuregs[16][26] ),
    .A1(_05725_),
    .S(_05897_),
    .X(_05900_));
 sky130_fd_sc_hd__clkbuf_1 _26255_ (.A(_05900_),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _26256_ (.A0(\cpuregs[16][27] ),
    .A1(_05727_),
    .S(_05897_),
    .X(_05901_));
 sky130_fd_sc_hd__clkbuf_1 _26257_ (.A(_05901_),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_1 _26258_ (.A0(\cpuregs[16][28] ),
    .A1(_05729_),
    .S(_05897_),
    .X(_05902_));
 sky130_fd_sc_hd__clkbuf_1 _26259_ (.A(_05902_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _26260_ (.A0(\cpuregs[16][29] ),
    .A1(_05731_),
    .S(_05897_),
    .X(_05903_));
 sky130_fd_sc_hd__clkbuf_1 _26261_ (.A(_05903_),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _26262_ (.A0(\cpuregs[16][30] ),
    .A1(_05733_),
    .S(_05868_),
    .X(_05904_));
 sky130_fd_sc_hd__clkbuf_1 _26263_ (.A(_05904_),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _26264_ (.A0(\cpuregs[16][31] ),
    .A1(_05735_),
    .S(_05868_),
    .X(_05905_));
 sky130_fd_sc_hd__clkbuf_1 _26265_ (.A(_05905_),
    .X(_00580_));
 sky130_fd_sc_hd__nor2_1 _26266_ (.A(_05340_),
    .B(_05866_),
    .Y(_05906_));
 sky130_fd_sc_hd__clkbuf_2 _26267_ (.A(_05906_),
    .X(_05907_));
 sky130_fd_sc_hd__buf_2 _26268_ (.A(_05907_),
    .X(_05908_));
 sky130_fd_sc_hd__mux2_1 _26269_ (.A0(\cpuregs[17][0] ),
    .A1(_05665_),
    .S(_05908_),
    .X(_05909_));
 sky130_fd_sc_hd__clkbuf_1 _26270_ (.A(_05909_),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _26271_ (.A0(\cpuregs[17][1] ),
    .A1(_05671_),
    .S(_05908_),
    .X(_05910_));
 sky130_fd_sc_hd__clkbuf_1 _26272_ (.A(_05910_),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _26273_ (.A0(\cpuregs[17][2] ),
    .A1(_05673_),
    .S(_05908_),
    .X(_05911_));
 sky130_fd_sc_hd__clkbuf_1 _26274_ (.A(_05911_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _26275_ (.A0(\cpuregs[17][3] ),
    .A1(_05675_),
    .S(_05908_),
    .X(_05912_));
 sky130_fd_sc_hd__clkbuf_1 _26276_ (.A(_05912_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _26277_ (.A0(\cpuregs[17][4] ),
    .A1(_05677_),
    .S(_05908_),
    .X(_05913_));
 sky130_fd_sc_hd__clkbuf_1 _26278_ (.A(_05913_),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _26279_ (.A0(\cpuregs[17][5] ),
    .A1(_05679_),
    .S(_05908_),
    .X(_05914_));
 sky130_fd_sc_hd__clkbuf_1 _26280_ (.A(_05914_),
    .X(_00586_));
 sky130_fd_sc_hd__buf_2 _26281_ (.A(_05907_),
    .X(_05915_));
 sky130_fd_sc_hd__mux2_1 _26282_ (.A0(\cpuregs[17][6] ),
    .A1(_05681_),
    .S(_05915_),
    .X(_05916_));
 sky130_fd_sc_hd__clkbuf_1 _26283_ (.A(_05916_),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _26284_ (.A0(\cpuregs[17][7] ),
    .A1(_05684_),
    .S(_05915_),
    .X(_05917_));
 sky130_fd_sc_hd__clkbuf_1 _26285_ (.A(_05917_),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _26286_ (.A0(\cpuregs[17][8] ),
    .A1(_05686_),
    .S(_05915_),
    .X(_05918_));
 sky130_fd_sc_hd__clkbuf_1 _26287_ (.A(_05918_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _26288_ (.A0(\cpuregs[17][9] ),
    .A1(_05688_),
    .S(_05915_),
    .X(_05919_));
 sky130_fd_sc_hd__clkbuf_1 _26289_ (.A(_05919_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _26290_ (.A0(\cpuregs[17][10] ),
    .A1(_05690_),
    .S(_05915_),
    .X(_05920_));
 sky130_fd_sc_hd__clkbuf_1 _26291_ (.A(_05920_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _26292_ (.A0(\cpuregs[17][11] ),
    .A1(_05692_),
    .S(_05915_),
    .X(_05921_));
 sky130_fd_sc_hd__clkbuf_1 _26293_ (.A(_05921_),
    .X(_00592_));
 sky130_fd_sc_hd__buf_2 _26294_ (.A(_05907_),
    .X(_05922_));
 sky130_fd_sc_hd__mux2_1 _26295_ (.A0(\cpuregs[17][12] ),
    .A1(_05694_),
    .S(_05922_),
    .X(_05923_));
 sky130_fd_sc_hd__clkbuf_1 _26296_ (.A(_05923_),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _26297_ (.A0(\cpuregs[17][13] ),
    .A1(_05697_),
    .S(_05922_),
    .X(_05924_));
 sky130_fd_sc_hd__clkbuf_1 _26298_ (.A(_05924_),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _26299_ (.A0(\cpuregs[17][14] ),
    .A1(_05699_),
    .S(_05922_),
    .X(_05925_));
 sky130_fd_sc_hd__clkbuf_1 _26300_ (.A(_05925_),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _26301_ (.A0(\cpuregs[17][15] ),
    .A1(_05701_),
    .S(_05922_),
    .X(_05926_));
 sky130_fd_sc_hd__clkbuf_1 _26302_ (.A(_05926_),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _26303_ (.A0(\cpuregs[17][16] ),
    .A1(_05703_),
    .S(_05922_),
    .X(_05927_));
 sky130_fd_sc_hd__clkbuf_1 _26304_ (.A(_05927_),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _26305_ (.A0(\cpuregs[17][17] ),
    .A1(_05705_),
    .S(_05922_),
    .X(_05928_));
 sky130_fd_sc_hd__clkbuf_1 _26306_ (.A(_05928_),
    .X(_00598_));
 sky130_fd_sc_hd__buf_2 _26307_ (.A(_05907_),
    .X(_05929_));
 sky130_fd_sc_hd__mux2_1 _26308_ (.A0(\cpuregs[17][18] ),
    .A1(_05707_),
    .S(_05929_),
    .X(_05930_));
 sky130_fd_sc_hd__clkbuf_1 _26309_ (.A(_05930_),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _26310_ (.A0(\cpuregs[17][19] ),
    .A1(_05710_),
    .S(_05929_),
    .X(_05931_));
 sky130_fd_sc_hd__clkbuf_1 _26311_ (.A(_05931_),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _26312_ (.A0(\cpuregs[17][20] ),
    .A1(_05712_),
    .S(_05929_),
    .X(_05932_));
 sky130_fd_sc_hd__clkbuf_1 _26313_ (.A(_05932_),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _26314_ (.A0(\cpuregs[17][21] ),
    .A1(_05714_),
    .S(_05929_),
    .X(_05933_));
 sky130_fd_sc_hd__clkbuf_1 _26315_ (.A(_05933_),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _26316_ (.A0(\cpuregs[17][22] ),
    .A1(_05716_),
    .S(_05929_),
    .X(_05934_));
 sky130_fd_sc_hd__clkbuf_1 _26317_ (.A(_05934_),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _26318_ (.A0(\cpuregs[17][23] ),
    .A1(_05718_),
    .S(_05929_),
    .X(_05935_));
 sky130_fd_sc_hd__clkbuf_1 _26319_ (.A(_05935_),
    .X(_00604_));
 sky130_fd_sc_hd__buf_2 _26320_ (.A(_05906_),
    .X(_05936_));
 sky130_fd_sc_hd__mux2_1 _26321_ (.A0(\cpuregs[17][24] ),
    .A1(_05720_),
    .S(_05936_),
    .X(_05937_));
 sky130_fd_sc_hd__clkbuf_1 _26322_ (.A(_05937_),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_1 _26323_ (.A0(\cpuregs[17][25] ),
    .A1(_05723_),
    .S(_05936_),
    .X(_05938_));
 sky130_fd_sc_hd__clkbuf_1 _26324_ (.A(_05938_),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_1 _26325_ (.A0(\cpuregs[17][26] ),
    .A1(_05725_),
    .S(_05936_),
    .X(_05939_));
 sky130_fd_sc_hd__clkbuf_1 _26326_ (.A(_05939_),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _26327_ (.A0(\cpuregs[17][27] ),
    .A1(_05727_),
    .S(_05936_),
    .X(_05940_));
 sky130_fd_sc_hd__clkbuf_1 _26328_ (.A(_05940_),
    .X(_00608_));
 sky130_fd_sc_hd__mux2_1 _26329_ (.A0(\cpuregs[17][28] ),
    .A1(_05729_),
    .S(_05936_),
    .X(_05941_));
 sky130_fd_sc_hd__clkbuf_1 _26330_ (.A(_05941_),
    .X(_00609_));
 sky130_fd_sc_hd__mux2_1 _26331_ (.A0(\cpuregs[17][29] ),
    .A1(_05731_),
    .S(_05936_),
    .X(_05942_));
 sky130_fd_sc_hd__clkbuf_1 _26332_ (.A(_05942_),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_1 _26333_ (.A0(\cpuregs[17][30] ),
    .A1(_05733_),
    .S(_05907_),
    .X(_05943_));
 sky130_fd_sc_hd__clkbuf_1 _26334_ (.A(_05943_),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _26335_ (.A0(\cpuregs[17][31] ),
    .A1(_05735_),
    .S(_05907_),
    .X(_05944_));
 sky130_fd_sc_hd__clkbuf_1 _26336_ (.A(_05944_),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_1 _26337_ (.A0(net33),
    .A1(\mem_rdata_q[0] ),
    .S(_05508_),
    .X(_05945_));
 sky130_fd_sc_hd__buf_1 _26338_ (.A(_05945_),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_1 _26339_ (.A0(net44),
    .A1(\mem_rdata_q[1] ),
    .S(_05508_),
    .X(_05946_));
 sky130_fd_sc_hd__clkbuf_1 _26340_ (.A(_05946_),
    .X(_00614_));
 sky130_fd_sc_hd__mux2_1 _26341_ (.A0(net55),
    .A1(\mem_rdata_q[2] ),
    .S(_05508_),
    .X(_05947_));
 sky130_fd_sc_hd__clkbuf_1 _26342_ (.A(_05947_),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _26343_ (.A0(net58),
    .A1(\mem_rdata_q[3] ),
    .S(_05523_),
    .X(_05948_));
 sky130_fd_sc_hd__buf_1 _26344_ (.A(_05948_),
    .X(_00616_));
 sky130_fd_sc_hd__mux2_1 _26345_ (.A0(net59),
    .A1(\mem_rdata_q[4] ),
    .S(_05523_),
    .X(_05949_));
 sky130_fd_sc_hd__buf_1 _26346_ (.A(_05949_),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _26347_ (.A0(net60),
    .A1(\mem_rdata_q[5] ),
    .S(_05523_),
    .X(_05950_));
 sky130_fd_sc_hd__buf_1 _26348_ (.A(_05950_),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _26349_ (.A0(net61),
    .A1(\mem_rdata_q[6] ),
    .S(_05523_),
    .X(_05951_));
 sky130_fd_sc_hd__buf_1 _26350_ (.A(_05951_),
    .X(_00619_));
 sky130_fd_sc_hd__clkbuf_2 _26351_ (.A(_05509_),
    .X(_05952_));
 sky130_fd_sc_hd__mux2_1 _26352_ (.A0(net62),
    .A1(\mem_rdata_q[7] ),
    .S(_05952_),
    .X(_05953_));
 sky130_fd_sc_hd__clkbuf_2 _26353_ (.A(_05953_),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _26354_ (.A0(net63),
    .A1(\mem_rdata_q[8] ),
    .S(_05952_),
    .X(_05954_));
 sky130_fd_sc_hd__clkbuf_2 _26355_ (.A(_05954_),
    .X(_00621_));
 sky130_fd_sc_hd__mux2_1 _26356_ (.A0(net64),
    .A1(\mem_rdata_q[9] ),
    .S(_05952_),
    .X(_05955_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26357_ (.A(_05955_),
    .X(_00622_));
 sky130_fd_sc_hd__mux2_1 _26358_ (.A0(net34),
    .A1(\mem_rdata_q[10] ),
    .S(_05952_),
    .X(_05956_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26359_ (.A(_05956_),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _26360_ (.A0(net35),
    .A1(\mem_rdata_q[11] ),
    .S(_05952_),
    .X(_05957_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26361_ (.A(_05957_),
    .X(_00624_));
 sky130_fd_sc_hd__mux2_1 _26362_ (.A0(net45),
    .A1(\mem_rdata_q[20] ),
    .S(_05952_),
    .X(_05958_));
 sky130_fd_sc_hd__clkbuf_1 _26363_ (.A(_05958_),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _26364_ (.A0(net46),
    .A1(\mem_rdata_q[21] ),
    .S(_05529_),
    .X(_05959_));
 sky130_fd_sc_hd__clkbuf_1 _26365_ (.A(_05959_),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _26366_ (.A0(net47),
    .A1(\mem_rdata_q[22] ),
    .S(_05529_),
    .X(_05960_));
 sky130_fd_sc_hd__clkbuf_1 _26367_ (.A(_05960_),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _26368_ (.A0(net48),
    .A1(\mem_rdata_q[23] ),
    .S(_05529_),
    .X(_05961_));
 sky130_fd_sc_hd__clkbuf_1 _26369_ (.A(_05961_),
    .X(_00636_));
 sky130_fd_sc_hd__nor2_1 _26370_ (.A(_05381_),
    .B(_05866_),
    .Y(_05962_));
 sky130_fd_sc_hd__buf_2 _26371_ (.A(_05962_),
    .X(_05963_));
 sky130_fd_sc_hd__buf_2 _26372_ (.A(_05963_),
    .X(_05964_));
 sky130_fd_sc_hd__mux2_1 _26373_ (.A0(\cpuregs[18][0] ),
    .A1(_05665_),
    .S(_05964_),
    .X(_05965_));
 sky130_fd_sc_hd__clkbuf_1 _26374_ (.A(_05965_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _26375_ (.A0(\cpuregs[18][1] ),
    .A1(_05671_),
    .S(_05964_),
    .X(_05966_));
 sky130_fd_sc_hd__clkbuf_1 _26376_ (.A(_05966_),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_1 _26377_ (.A0(\cpuregs[18][2] ),
    .A1(_05673_),
    .S(_05964_),
    .X(_05967_));
 sky130_fd_sc_hd__clkbuf_1 _26378_ (.A(_05967_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _26379_ (.A0(\cpuregs[18][3] ),
    .A1(_05675_),
    .S(_05964_),
    .X(_05968_));
 sky130_fd_sc_hd__clkbuf_1 _26380_ (.A(_05968_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _26381_ (.A0(\cpuregs[18][4] ),
    .A1(_05677_),
    .S(_05964_),
    .X(_05969_));
 sky130_fd_sc_hd__clkbuf_1 _26382_ (.A(_05969_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _26383_ (.A0(\cpuregs[18][5] ),
    .A1(_05679_),
    .S(_05964_),
    .X(_05970_));
 sky130_fd_sc_hd__clkbuf_1 _26384_ (.A(_05970_),
    .X(_00650_));
 sky130_fd_sc_hd__buf_2 _26385_ (.A(_05963_),
    .X(_05971_));
 sky130_fd_sc_hd__mux2_1 _26386_ (.A0(\cpuregs[18][6] ),
    .A1(_05681_),
    .S(_05971_),
    .X(_05972_));
 sky130_fd_sc_hd__clkbuf_1 _26387_ (.A(_05972_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _26388_ (.A0(\cpuregs[18][7] ),
    .A1(_05684_),
    .S(_05971_),
    .X(_05973_));
 sky130_fd_sc_hd__clkbuf_1 _26389_ (.A(_05973_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _26390_ (.A0(\cpuregs[18][8] ),
    .A1(_05686_),
    .S(_05971_),
    .X(_05974_));
 sky130_fd_sc_hd__clkbuf_1 _26391_ (.A(_05974_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _26392_ (.A0(\cpuregs[18][9] ),
    .A1(_05688_),
    .S(_05971_),
    .X(_05975_));
 sky130_fd_sc_hd__clkbuf_1 _26393_ (.A(_05975_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _26394_ (.A0(\cpuregs[18][10] ),
    .A1(_05690_),
    .S(_05971_),
    .X(_05976_));
 sky130_fd_sc_hd__clkbuf_1 _26395_ (.A(_05976_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _26396_ (.A0(\cpuregs[18][11] ),
    .A1(_05692_),
    .S(_05971_),
    .X(_05977_));
 sky130_fd_sc_hd__clkbuf_1 _26397_ (.A(_05977_),
    .X(_00656_));
 sky130_fd_sc_hd__buf_2 _26398_ (.A(_05963_),
    .X(_05978_));
 sky130_fd_sc_hd__mux2_1 _26399_ (.A0(\cpuregs[18][12] ),
    .A1(_05694_),
    .S(_05978_),
    .X(_05979_));
 sky130_fd_sc_hd__clkbuf_1 _26400_ (.A(_05979_),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _26401_ (.A0(\cpuregs[18][13] ),
    .A1(_05697_),
    .S(_05978_),
    .X(_05980_));
 sky130_fd_sc_hd__clkbuf_1 _26402_ (.A(_05980_),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _26403_ (.A0(\cpuregs[18][14] ),
    .A1(_05699_),
    .S(_05978_),
    .X(_05981_));
 sky130_fd_sc_hd__clkbuf_1 _26404_ (.A(_05981_),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _26405_ (.A0(\cpuregs[18][15] ),
    .A1(_05701_),
    .S(_05978_),
    .X(_05982_));
 sky130_fd_sc_hd__clkbuf_1 _26406_ (.A(_05982_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _26407_ (.A0(\cpuregs[18][16] ),
    .A1(_05703_),
    .S(_05978_),
    .X(_05983_));
 sky130_fd_sc_hd__clkbuf_1 _26408_ (.A(_05983_),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _26409_ (.A0(\cpuregs[18][17] ),
    .A1(_05705_),
    .S(_05978_),
    .X(_05984_));
 sky130_fd_sc_hd__clkbuf_1 _26410_ (.A(_05984_),
    .X(_00662_));
 sky130_fd_sc_hd__buf_2 _26411_ (.A(_05963_),
    .X(_05985_));
 sky130_fd_sc_hd__mux2_1 _26412_ (.A0(\cpuregs[18][18] ),
    .A1(_05707_),
    .S(_05985_),
    .X(_05986_));
 sky130_fd_sc_hd__clkbuf_1 _26413_ (.A(_05986_),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _26414_ (.A0(\cpuregs[18][19] ),
    .A1(_05710_),
    .S(_05985_),
    .X(_05987_));
 sky130_fd_sc_hd__clkbuf_1 _26415_ (.A(_05987_),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _26416_ (.A0(\cpuregs[18][20] ),
    .A1(_05712_),
    .S(_05985_),
    .X(_05988_));
 sky130_fd_sc_hd__clkbuf_1 _26417_ (.A(_05988_),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_1 _26418_ (.A0(\cpuregs[18][21] ),
    .A1(_05714_),
    .S(_05985_),
    .X(_05989_));
 sky130_fd_sc_hd__clkbuf_1 _26419_ (.A(_05989_),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_1 _26420_ (.A0(\cpuregs[18][22] ),
    .A1(_05716_),
    .S(_05985_),
    .X(_05990_));
 sky130_fd_sc_hd__clkbuf_1 _26421_ (.A(_05990_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _26422_ (.A0(\cpuregs[18][23] ),
    .A1(_05718_),
    .S(_05985_),
    .X(_05991_));
 sky130_fd_sc_hd__clkbuf_1 _26423_ (.A(_05991_),
    .X(_00668_));
 sky130_fd_sc_hd__buf_2 _26424_ (.A(_05962_),
    .X(_05992_));
 sky130_fd_sc_hd__mux2_1 _26425_ (.A0(\cpuregs[18][24] ),
    .A1(_05720_),
    .S(_05992_),
    .X(_05993_));
 sky130_fd_sc_hd__clkbuf_1 _26426_ (.A(_05993_),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _26427_ (.A0(\cpuregs[18][25] ),
    .A1(_05723_),
    .S(_05992_),
    .X(_05994_));
 sky130_fd_sc_hd__clkbuf_1 _26428_ (.A(_05994_),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_1 _26429_ (.A0(\cpuregs[18][26] ),
    .A1(_05725_),
    .S(_05992_),
    .X(_05995_));
 sky130_fd_sc_hd__clkbuf_1 _26430_ (.A(_05995_),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_1 _26431_ (.A0(\cpuregs[18][27] ),
    .A1(_05727_),
    .S(_05992_),
    .X(_05996_));
 sky130_fd_sc_hd__clkbuf_1 _26432_ (.A(_05996_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _26433_ (.A0(\cpuregs[18][28] ),
    .A1(_05729_),
    .S(_05992_),
    .X(_05997_));
 sky130_fd_sc_hd__clkbuf_1 _26434_ (.A(_05997_),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _26435_ (.A0(\cpuregs[18][29] ),
    .A1(_05731_),
    .S(_05992_),
    .X(_05998_));
 sky130_fd_sc_hd__clkbuf_1 _26436_ (.A(_05998_),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _26437_ (.A0(\cpuregs[18][30] ),
    .A1(_05733_),
    .S(_05963_),
    .X(_05999_));
 sky130_fd_sc_hd__clkbuf_1 _26438_ (.A(_05999_),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _26439_ (.A0(\cpuregs[18][31] ),
    .A1(_05735_),
    .S(_05963_),
    .X(_06000_));
 sky130_fd_sc_hd__clkbuf_1 _26440_ (.A(_06000_),
    .X(_00676_));
 sky130_fd_sc_hd__nor2_1 _26441_ (.A(_05269_),
    .B(_05381_),
    .Y(_06001_));
 sky130_fd_sc_hd__buf_4 _26442_ (.A(_06001_),
    .X(_06002_));
 sky130_fd_sc_hd__buf_2 _26443_ (.A(_06002_),
    .X(_06003_));
 sky130_fd_sc_hd__mux2_1 _26444_ (.A0(\cpuregs[2][0] ),
    .A1(_05665_),
    .S(_06003_),
    .X(_06004_));
 sky130_fd_sc_hd__clkbuf_1 _26445_ (.A(_06004_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _26446_ (.A0(\cpuregs[2][1] ),
    .A1(_05671_),
    .S(_06003_),
    .X(_06005_));
 sky130_fd_sc_hd__clkbuf_1 _26447_ (.A(_06005_),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _26448_ (.A0(\cpuregs[2][2] ),
    .A1(_05673_),
    .S(_06003_),
    .X(_06006_));
 sky130_fd_sc_hd__clkbuf_1 _26449_ (.A(_06006_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _26450_ (.A0(\cpuregs[2][3] ),
    .A1(_05675_),
    .S(_06003_),
    .X(_06007_));
 sky130_fd_sc_hd__clkbuf_1 _26451_ (.A(_06007_),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _26452_ (.A0(\cpuregs[2][4] ),
    .A1(_05677_),
    .S(_06003_),
    .X(_06008_));
 sky130_fd_sc_hd__clkbuf_1 _26453_ (.A(_06008_),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _26454_ (.A0(\cpuregs[2][5] ),
    .A1(_05679_),
    .S(_06003_),
    .X(_06009_));
 sky130_fd_sc_hd__clkbuf_1 _26455_ (.A(_06009_),
    .X(_00682_));
 sky130_fd_sc_hd__clkbuf_4 _26456_ (.A(_06002_),
    .X(_06010_));
 sky130_fd_sc_hd__mux2_1 _26457_ (.A0(\cpuregs[2][6] ),
    .A1(_05681_),
    .S(_06010_),
    .X(_06011_));
 sky130_fd_sc_hd__clkbuf_1 _26458_ (.A(_06011_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _26459_ (.A0(\cpuregs[2][7] ),
    .A1(_05684_),
    .S(_06010_),
    .X(_06012_));
 sky130_fd_sc_hd__clkbuf_1 _26460_ (.A(_06012_),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _26461_ (.A0(\cpuregs[2][8] ),
    .A1(_05686_),
    .S(_06010_),
    .X(_06013_));
 sky130_fd_sc_hd__clkbuf_1 _26462_ (.A(_06013_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _26463_ (.A0(\cpuregs[2][9] ),
    .A1(_05688_),
    .S(_06010_),
    .X(_06014_));
 sky130_fd_sc_hd__clkbuf_1 _26464_ (.A(_06014_),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _26465_ (.A0(\cpuregs[2][10] ),
    .A1(_05690_),
    .S(_06010_),
    .X(_06015_));
 sky130_fd_sc_hd__clkbuf_1 _26466_ (.A(_06015_),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _26467_ (.A0(\cpuregs[2][11] ),
    .A1(_05692_),
    .S(_06010_),
    .X(_06016_));
 sky130_fd_sc_hd__clkbuf_1 _26468_ (.A(_06016_),
    .X(_00688_));
 sky130_fd_sc_hd__buf_2 _26469_ (.A(_06002_),
    .X(_06017_));
 sky130_fd_sc_hd__mux2_1 _26470_ (.A0(\cpuregs[2][12] ),
    .A1(_05694_),
    .S(_06017_),
    .X(_06018_));
 sky130_fd_sc_hd__clkbuf_1 _26471_ (.A(_06018_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _26472_ (.A0(\cpuregs[2][13] ),
    .A1(_05697_),
    .S(_06017_),
    .X(_06019_));
 sky130_fd_sc_hd__clkbuf_1 _26473_ (.A(_06019_),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _26474_ (.A0(\cpuregs[2][14] ),
    .A1(_05699_),
    .S(_06017_),
    .X(_06020_));
 sky130_fd_sc_hd__clkbuf_1 _26475_ (.A(_06020_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _26476_ (.A0(\cpuregs[2][15] ),
    .A1(_05701_),
    .S(_06017_),
    .X(_06021_));
 sky130_fd_sc_hd__clkbuf_1 _26477_ (.A(_06021_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _26478_ (.A0(\cpuregs[2][16] ),
    .A1(_05703_),
    .S(_06017_),
    .X(_06022_));
 sky130_fd_sc_hd__clkbuf_1 _26479_ (.A(_06022_),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _26480_ (.A0(\cpuregs[2][17] ),
    .A1(_05705_),
    .S(_06017_),
    .X(_06023_));
 sky130_fd_sc_hd__clkbuf_1 _26481_ (.A(_06023_),
    .X(_00694_));
 sky130_fd_sc_hd__buf_2 _26482_ (.A(_06002_),
    .X(_06024_));
 sky130_fd_sc_hd__mux2_1 _26483_ (.A0(\cpuregs[2][18] ),
    .A1(_05707_),
    .S(_06024_),
    .X(_06025_));
 sky130_fd_sc_hd__clkbuf_1 _26484_ (.A(_06025_),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _26485_ (.A0(\cpuregs[2][19] ),
    .A1(_05710_),
    .S(_06024_),
    .X(_06026_));
 sky130_fd_sc_hd__clkbuf_1 _26486_ (.A(_06026_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _26487_ (.A0(\cpuregs[2][20] ),
    .A1(_05712_),
    .S(_06024_),
    .X(_06027_));
 sky130_fd_sc_hd__clkbuf_1 _26488_ (.A(_06027_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _26489_ (.A0(\cpuregs[2][21] ),
    .A1(_05714_),
    .S(_06024_),
    .X(_06028_));
 sky130_fd_sc_hd__clkbuf_1 _26490_ (.A(_06028_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _26491_ (.A0(\cpuregs[2][22] ),
    .A1(_05716_),
    .S(_06024_),
    .X(_06029_));
 sky130_fd_sc_hd__clkbuf_1 _26492_ (.A(_06029_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _26493_ (.A0(\cpuregs[2][23] ),
    .A1(_05718_),
    .S(_06024_),
    .X(_06030_));
 sky130_fd_sc_hd__clkbuf_1 _26494_ (.A(_06030_),
    .X(_00700_));
 sky130_fd_sc_hd__clkbuf_4 _26495_ (.A(_06001_),
    .X(_06031_));
 sky130_fd_sc_hd__mux2_1 _26496_ (.A0(\cpuregs[2][24] ),
    .A1(_05720_),
    .S(_06031_),
    .X(_06032_));
 sky130_fd_sc_hd__clkbuf_1 _26497_ (.A(_06032_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _26498_ (.A0(\cpuregs[2][25] ),
    .A1(_05723_),
    .S(_06031_),
    .X(_06033_));
 sky130_fd_sc_hd__clkbuf_1 _26499_ (.A(_06033_),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_1 _26500_ (.A0(\cpuregs[2][26] ),
    .A1(_05725_),
    .S(_06031_),
    .X(_06034_));
 sky130_fd_sc_hd__clkbuf_1 _26501_ (.A(_06034_),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _26502_ (.A0(\cpuregs[2][27] ),
    .A1(_05727_),
    .S(_06031_),
    .X(_06035_));
 sky130_fd_sc_hd__clkbuf_1 _26503_ (.A(_06035_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _26504_ (.A0(\cpuregs[2][28] ),
    .A1(_05729_),
    .S(_06031_),
    .X(_06036_));
 sky130_fd_sc_hd__clkbuf_1 _26505_ (.A(_06036_),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _26506_ (.A0(\cpuregs[2][29] ),
    .A1(_05731_),
    .S(_06031_),
    .X(_06037_));
 sky130_fd_sc_hd__clkbuf_1 _26507_ (.A(_06037_),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _26508_ (.A0(\cpuregs[2][30] ),
    .A1(_05733_),
    .S(_06002_),
    .X(_06038_));
 sky130_fd_sc_hd__clkbuf_1 _26509_ (.A(_06038_),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _26510_ (.A0(\cpuregs[2][31] ),
    .A1(_05735_),
    .S(_06002_),
    .X(_06039_));
 sky130_fd_sc_hd__clkbuf_1 _26511_ (.A(_06039_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _26512_ (.A0(_10264_),
    .A1(_10603_),
    .S(_05425_),
    .X(_06040_));
 sky130_fd_sc_hd__clkbuf_1 _26513_ (.A(_06040_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _26514_ (.A0(_10104_),
    .A1(_10598_),
    .S(_05425_),
    .X(_06041_));
 sky130_fd_sc_hd__clkbuf_1 _26515_ (.A(_06041_),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _26516_ (.A0(_10311_),
    .A1(_10609_),
    .S(_05425_),
    .X(_06042_));
 sky130_fd_sc_hd__clkbuf_1 _26517_ (.A(_06042_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _26518_ (.A0(_10322_),
    .A1(_10651_),
    .S(_05425_),
    .X(_06043_));
 sky130_fd_sc_hd__clkbuf_1 _26519_ (.A(_06043_),
    .X(_00712_));
 sky130_fd_sc_hd__buf_2 _26520_ (.A(_05424_),
    .X(_06044_));
 sky130_fd_sc_hd__mux2_1 _26521_ (.A0(_10331_),
    .A1(_10667_),
    .S(_06044_),
    .X(_06045_));
 sky130_fd_sc_hd__clkbuf_1 _26522_ (.A(_06045_),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _26523_ (.A0(_10334_),
    .A1(_11343_),
    .S(_06044_),
    .X(_06046_));
 sky130_fd_sc_hd__clkbuf_1 _26524_ (.A(_06046_),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _26525_ (.A0(_10337_),
    .A1(_12361_),
    .S(_06044_),
    .X(_06047_));
 sky130_fd_sc_hd__clkbuf_1 _26526_ (.A(_06047_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _26527_ (.A0(_08461_),
    .A1(_11297_),
    .S(_06044_),
    .X(_06048_));
 sky130_fd_sc_hd__clkbuf_1 _26528_ (.A(_06048_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _26529_ (.A0(_10344_),
    .A1(_11050_),
    .S(_06044_),
    .X(_06049_));
 sky130_fd_sc_hd__clkbuf_1 _26530_ (.A(_06049_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _26531_ (.A0(_10157_),
    .A1(_11167_),
    .S(_06044_),
    .X(_06050_));
 sky130_fd_sc_hd__clkbuf_1 _26532_ (.A(_06050_),
    .X(_00718_));
 sky130_fd_sc_hd__clkbuf_2 _26533_ (.A(_05424_),
    .X(_06051_));
 sky130_fd_sc_hd__mux2_1 _26534_ (.A0(_10163_),
    .A1(_11157_),
    .S(_06051_),
    .X(_06052_));
 sky130_fd_sc_hd__clkbuf_1 _26535_ (.A(_06052_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _26536_ (.A0(_08412_),
    .A1(_11161_),
    .S(_06051_),
    .X(_06053_));
 sky130_fd_sc_hd__clkbuf_1 _26537_ (.A(_06053_),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _26538_ (.A0(_10354_),
    .A1(_11474_),
    .S(_06051_),
    .X(_06054_));
 sky130_fd_sc_hd__clkbuf_1 _26539_ (.A(_06054_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _26540_ (.A0(_10357_),
    .A1(_11369_),
    .S(_06051_),
    .X(_06055_));
 sky130_fd_sc_hd__clkbuf_1 _26541_ (.A(_06055_),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _26542_ (.A0(_10361_),
    .A1(_11382_),
    .S(_06051_),
    .X(_06056_));
 sky130_fd_sc_hd__clkbuf_1 _26543_ (.A(_06056_),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _26544_ (.A0(_10187_),
    .A1(_11826_),
    .S(_06051_),
    .X(_06057_));
 sky130_fd_sc_hd__clkbuf_1 _26545_ (.A(_06057_),
    .X(_00724_));
 sky130_fd_sc_hd__clkbuf_4 _26546_ (.A(_05424_),
    .X(_06058_));
 sky130_fd_sc_hd__mux2_1 _26547_ (.A0(_10367_),
    .A1(_11954_),
    .S(_06058_),
    .X(_06059_));
 sky130_fd_sc_hd__buf_1 _26548_ (.A(_06059_),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _26549_ (.A0(_10197_),
    .A1(_13919_),
    .S(_06058_),
    .X(_06060_));
 sky130_fd_sc_hd__buf_1 _26550_ (.A(_06060_),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _26551_ (.A0(_10372_),
    .A1(_14283_),
    .S(_06058_),
    .X(_06061_));
 sky130_fd_sc_hd__buf_1 _26552_ (.A(_06061_),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _26553_ (.A0(_10206_),
    .A1(_14457_),
    .S(_06058_),
    .X(_06062_));
 sky130_fd_sc_hd__clkbuf_2 _26554_ (.A(_06062_),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _26555_ (.A0(_10378_),
    .A1(_01558_),
    .S(_06058_),
    .X(_06063_));
 sky130_fd_sc_hd__clkbuf_1 _26556_ (.A(_06063_),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _26557_ (.A0(_10214_),
    .A1(_01564_),
    .S(_06058_),
    .X(_06064_));
 sky130_fd_sc_hd__clkbuf_1 _26558_ (.A(_06064_),
    .X(_00730_));
 sky130_fd_sc_hd__buf_2 _26559_ (.A(_05424_),
    .X(_06065_));
 sky130_fd_sc_hd__mux2_1 _26560_ (.A0(_10384_),
    .A1(_01885_),
    .S(_06065_),
    .X(_06066_));
 sky130_fd_sc_hd__clkbuf_1 _26561_ (.A(_06066_),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _26562_ (.A0(_10224_),
    .A1(_02036_),
    .S(_06065_),
    .X(_06067_));
 sky130_fd_sc_hd__clkbuf_1 _26563_ (.A(_06067_),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _26564_ (.A0(_10389_),
    .A1(_03308_),
    .S(_06065_),
    .X(_06068_));
 sky130_fd_sc_hd__clkbuf_1 _26565_ (.A(_06068_),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _26566_ (.A0(_10392_),
    .A1(_02331_),
    .S(_06065_),
    .X(_06069_));
 sky130_fd_sc_hd__clkbuf_1 _26567_ (.A(_06069_),
    .X(_00734_));
 sky130_fd_sc_hd__mux2_1 _26568_ (.A0(_10397_),
    .A1(_02472_),
    .S(_06065_),
    .X(_06070_));
 sky130_fd_sc_hd__clkbuf_1 _26569_ (.A(_06070_),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_1 _26570_ (.A0(_10241_),
    .A1(_04092_),
    .S(_06065_),
    .X(_06071_));
 sky130_fd_sc_hd__clkbuf_1 _26571_ (.A(_06071_),
    .X(_00736_));
 sky130_fd_sc_hd__buf_2 _26572_ (.A(_05424_),
    .X(_06072_));
 sky130_fd_sc_hd__mux2_1 _26573_ (.A0(_10246_),
    .A1(_04090_),
    .S(_06072_),
    .X(_06073_));
 sky130_fd_sc_hd__clkbuf_1 _26574_ (.A(_06073_),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_1 _26575_ (.A0(_10250_),
    .A1(_13816_),
    .S(_06072_),
    .X(_06074_));
 sky130_fd_sc_hd__buf_1 _26576_ (.A(_06074_),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_1 _26577_ (.A0(_10255_),
    .A1(_13819_),
    .S(_06072_),
    .X(_06075_));
 sky130_fd_sc_hd__clkbuf_1 _26578_ (.A(_06075_),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_1 _26579_ (.A0(_10259_),
    .A1(_14214_),
    .S(_06072_),
    .X(_06076_));
 sky130_fd_sc_hd__clkbuf_1 _26580_ (.A(_06076_),
    .X(_00740_));
 sky130_fd_sc_hd__mux2_1 _26581_ (.A0(_10270_),
    .A1(_10586_),
    .S(_06072_),
    .X(_06077_));
 sky130_fd_sc_hd__clkbuf_1 _26582_ (.A(_06077_),
    .X(_00741_));
 sky130_fd_sc_hd__mux2_1 _26583_ (.A0(_10108_),
    .A1(_10602_),
    .S(_06072_),
    .X(_06078_));
 sky130_fd_sc_hd__clkbuf_1 _26584_ (.A(_06078_),
    .X(_00742_));
 sky130_fd_sc_hd__clkbuf_2 _26585_ (.A(_05423_),
    .X(_06079_));
 sky130_fd_sc_hd__mux2_1 _26586_ (.A0(_10273_),
    .A1(_10613_),
    .S(_06079_),
    .X(_06080_));
 sky130_fd_sc_hd__clkbuf_1 _26587_ (.A(_06080_),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_1 _26588_ (.A0(_04961_),
    .A1(_11368_),
    .S(_06079_),
    .X(_06081_));
 sky130_fd_sc_hd__clkbuf_1 _26589_ (.A(_06081_),
    .X(_00744_));
 sky130_fd_sc_hd__mux2_1 _26590_ (.A0(_04755_),
    .A1(_10663_),
    .S(_06079_),
    .X(_06082_));
 sky130_fd_sc_hd__clkbuf_1 _26591_ (.A(_06082_),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_1 _26592_ (.A0(_10277_),
    .A1(_14223_),
    .S(_06079_),
    .X(_06083_));
 sky130_fd_sc_hd__clkbuf_1 _26593_ (.A(_06083_),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _26594_ (.A0(_10279_),
    .A1(_10738_),
    .S(_06079_),
    .X(_06084_));
 sky130_fd_sc_hd__clkbuf_1 _26595_ (.A(_06084_),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _26596_ (.A0(_10280_),
    .A1(_10784_),
    .S(_06079_),
    .X(_06085_));
 sky130_fd_sc_hd__clkbuf_1 _26597_ (.A(_06085_),
    .X(_00748_));
 sky130_fd_sc_hd__buf_2 _26598_ (.A(_05423_),
    .X(_06086_));
 sky130_fd_sc_hd__mux2_1 _26599_ (.A0(_08484_),
    .A1(_13858_),
    .S(_06086_),
    .X(_06087_));
 sky130_fd_sc_hd__clkbuf_1 _26600_ (.A(_06087_),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _26601_ (.A0(_10158_),
    .A1(_10895_),
    .S(_06086_),
    .X(_06088_));
 sky130_fd_sc_hd__clkbuf_1 _26602_ (.A(_06088_),
    .X(_00750_));
 sky130_fd_sc_hd__mux2_1 _26603_ (.A0(_10164_),
    .A1(_10958_),
    .S(_06086_),
    .X(_06089_));
 sky130_fd_sc_hd__clkbuf_1 _26604_ (.A(_06089_),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_1 _26605_ (.A0(_08413_),
    .A1(_11109_),
    .S(_06086_),
    .X(_06090_));
 sky130_fd_sc_hd__clkbuf_1 _26606_ (.A(_06090_),
    .X(_00752_));
 sky130_fd_sc_hd__mux2_1 _26607_ (.A0(_08343_),
    .A1(_11137_),
    .S(_06086_),
    .X(_06091_));
 sky130_fd_sc_hd__clkbuf_1 _26608_ (.A(_06091_),
    .X(_00753_));
 sky130_fd_sc_hd__mux2_1 _26609_ (.A0(_08347_),
    .A1(_11237_),
    .S(_06086_),
    .X(_06092_));
 sky130_fd_sc_hd__clkbuf_1 _26610_ (.A(_06092_),
    .X(_00754_));
 sky130_fd_sc_hd__clkbuf_2 _26611_ (.A(_05423_),
    .X(_06093_));
 sky130_fd_sc_hd__mux2_1 _26612_ (.A0(_08419_),
    .A1(_01547_),
    .S(_06093_),
    .X(_06094_));
 sky130_fd_sc_hd__clkbuf_1 _26613_ (.A(_06094_),
    .X(_00755_));
 sky130_fd_sc_hd__mux2_1 _26614_ (.A0(_10188_),
    .A1(_11447_),
    .S(_06093_),
    .X(_06095_));
 sky130_fd_sc_hd__clkbuf_1 _26615_ (.A(_06095_),
    .X(_00756_));
 sky130_fd_sc_hd__mux2_1 _26616_ (.A0(net306),
    .A1(_11557_),
    .S(_06093_),
    .X(_06096_));
 sky130_fd_sc_hd__clkbuf_1 _26617_ (.A(_06096_),
    .X(_00757_));
 sky130_fd_sc_hd__mux2_1 _26618_ (.A0(_08383_),
    .A1(_11666_),
    .S(_06093_),
    .X(_06097_));
 sky130_fd_sc_hd__clkbuf_1 _26619_ (.A(_06097_),
    .X(_00758_));
 sky130_fd_sc_hd__mux2_1 _26620_ (.A0(net308),
    .A1(_11773_),
    .S(_06093_),
    .X(_06098_));
 sky130_fd_sc_hd__clkbuf_1 _26621_ (.A(_06098_),
    .X(_00759_));
 sky130_fd_sc_hd__mux2_1 _26622_ (.A0(_08375_),
    .A1(_11892_),
    .S(_06093_),
    .X(_06099_));
 sky130_fd_sc_hd__clkbuf_1 _26623_ (.A(_06099_),
    .X(_00760_));
 sky130_fd_sc_hd__buf_2 _26624_ (.A(_05423_),
    .X(_06100_));
 sky130_fd_sc_hd__mux2_1 _26625_ (.A0(net311),
    .A1(_01583_),
    .S(_06100_),
    .X(_06101_));
 sky130_fd_sc_hd__clkbuf_1 _26626_ (.A(_06101_),
    .X(_00761_));
 sky130_fd_sc_hd__mux2_1 _26627_ (.A0(_08364_),
    .A1(_12229_),
    .S(_06100_),
    .X(_06102_));
 sky130_fd_sc_hd__clkbuf_1 _26628_ (.A(_06102_),
    .X(_00762_));
 sky130_fd_sc_hd__mux2_1 _26629_ (.A0(net313),
    .A1(_12325_),
    .S(_06100_),
    .X(_06103_));
 sky130_fd_sc_hd__clkbuf_1 _26630_ (.A(_06103_),
    .X(_00763_));
 sky130_fd_sc_hd__mux2_1 _26631_ (.A0(_08369_),
    .A1(_03633_),
    .S(_06100_),
    .X(_06104_));
 sky130_fd_sc_hd__clkbuf_1 _26632_ (.A(_06104_),
    .X(_00764_));
 sky130_fd_sc_hd__mux2_1 _26633_ (.A0(net315),
    .A1(_12587_),
    .S(_06100_),
    .X(_06105_));
 sky130_fd_sc_hd__clkbuf_1 _26634_ (.A(_06105_),
    .X(_00765_));
 sky130_fd_sc_hd__mux2_1 _26635_ (.A0(_08427_),
    .A1(_12773_),
    .S(_06100_),
    .X(_06106_));
 sky130_fd_sc_hd__clkbuf_1 _26636_ (.A(_06106_),
    .X(_00766_));
 sky130_fd_sc_hd__clkbuf_2 _26637_ (.A(_05423_),
    .X(_06107_));
 sky130_fd_sc_hd__mux2_1 _26638_ (.A0(net317),
    .A1(_03609_),
    .S(_06107_),
    .X(_06108_));
 sky130_fd_sc_hd__buf_1 _26639_ (.A(_06108_),
    .X(_00767_));
 sky130_fd_sc_hd__mux2_2 _26640_ (.A0(_08436_),
    .A1(_04098_),
    .S(_06107_),
    .X(_06109_));
 sky130_fd_sc_hd__clkbuf_1 _26641_ (.A(_06109_),
    .X(_00768_));
 sky130_fd_sc_hd__mux2_2 _26642_ (.A0(_08479_),
    .A1(_04089_),
    .S(_06107_),
    .X(_06110_));
 sky130_fd_sc_hd__clkbuf_1 _26643_ (.A(_06110_),
    .X(_00769_));
 sky130_fd_sc_hd__mux2_2 _26644_ (.A0(_08398_),
    .A1(_04091_),
    .S(_06107_),
    .X(_06111_));
 sky130_fd_sc_hd__clkbuf_1 _26645_ (.A(_06111_),
    .X(_00770_));
 sky130_fd_sc_hd__mux2_1 _26646_ (.A0(_08487_),
    .A1(_04511_),
    .S(_06107_),
    .X(_06112_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26647_ (.A(_06112_),
    .X(_00771_));
 sky130_fd_sc_hd__mux2_2 _26648_ (.A0(_10260_),
    .A1(_04254_),
    .S(_06107_),
    .X(_06113_));
 sky130_fd_sc_hd__clkbuf_1 _26649_ (.A(_06113_),
    .X(_00772_));
 sky130_fd_sc_hd__clkbuf_4 _26650_ (.A(_08505_),
    .X(_06114_));
 sky130_fd_sc_hd__and2_1 _26651_ (.A(_06114_),
    .B(\genblk1.pcpi_mul.active[0] ),
    .X(_06115_));
 sky130_fd_sc_hd__clkbuf_1 _26652_ (.A(_06115_),
    .X(_00774_));
 sky130_fd_sc_hd__a21oi_1 _26653_ (.A1(net331),
    .A2(_08318_),
    .B1(_08516_),
    .Y(_06116_));
 sky130_fd_sc_hd__nor2_1 _26654_ (.A(_08521_),
    .B(_06116_),
    .Y(_00775_));
 sky130_fd_sc_hd__clkbuf_2 _26655_ (.A(_08145_),
    .X(_06117_));
 sky130_fd_sc_hd__or2_1 _26656_ (.A(\cpu_state[1] ),
    .B(\cpu_state[2] ),
    .X(_06118_));
 sky130_fd_sc_hd__or2_1 _26657_ (.A(_08513_),
    .B(instr_retirq),
    .X(_06119_));
 sky130_fd_sc_hd__o211a_1 _26658_ (.A1(_04977_),
    .A2(_06117_),
    .B1(_06118_),
    .C1(_06119_),
    .X(_06120_));
 sky130_fd_sc_hd__buf_1 _26659_ (.A(_06120_),
    .X(_06121_));
 sky130_fd_sc_hd__clkbuf_2 _26660_ (.A(_06121_),
    .X(_06122_));
 sky130_fd_sc_hd__clkbuf_2 _26661_ (.A(_06122_),
    .X(_06123_));
 sky130_fd_sc_hd__clkbuf_2 _26662_ (.A(_08513_),
    .X(_06124_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26663_ (.A(_06124_),
    .X(_06125_));
 sky130_fd_sc_hd__clkbuf_2 _26664_ (.A(_06125_),
    .X(_06126_));
 sky130_fd_sc_hd__buf_1 _26665_ (.A(_06120_),
    .X(_06127_));
 sky130_fd_sc_hd__a21bo_1 _26666_ (.A1(_06126_),
    .A2(_08240_),
    .B1_N(_06127_),
    .X(_06128_));
 sky130_fd_sc_hd__buf_2 _26667_ (.A(_08505_),
    .X(_06129_));
 sky130_fd_sc_hd__buf_2 _26668_ (.A(_06129_),
    .X(_06130_));
 sky130_fd_sc_hd__o211a_1 _26669_ (.A1(net67),
    .A2(_06123_),
    .B1(_06128_),
    .C1(_06130_),
    .X(_00776_));
 sky130_fd_sc_hd__a21bo_1 _26670_ (.A1(_06126_),
    .A2(_08263_),
    .B1_N(_06127_),
    .X(_06131_));
 sky130_fd_sc_hd__o211a_1 _26671_ (.A1(net78),
    .A2(_06123_),
    .B1(_06131_),
    .C1(_06130_),
    .X(_00777_));
 sky130_fd_sc_hd__a21bo_1 _26672_ (.A1(_06126_),
    .A2(_08268_),
    .B1_N(_06127_),
    .X(_06132_));
 sky130_fd_sc_hd__o211a_1 _26673_ (.A1(net89),
    .A2(_06123_),
    .B1(_06132_),
    .C1(_06130_),
    .X(_00778_));
 sky130_fd_sc_hd__a21bo_1 _26674_ (.A1(_06126_),
    .A2(_08236_),
    .B1_N(_06127_),
    .X(_06133_));
 sky130_fd_sc_hd__o211a_1 _26675_ (.A1(net92),
    .A2(_06123_),
    .B1(_06133_),
    .C1(_06130_),
    .X(_00779_));
 sky130_fd_sc_hd__a21bo_1 _26676_ (.A1(_06126_),
    .A2(_08267_),
    .B1_N(_06127_),
    .X(_06134_));
 sky130_fd_sc_hd__clkbuf_2 _26677_ (.A(_06114_),
    .X(_06135_));
 sky130_fd_sc_hd__o211a_1 _26678_ (.A1(net93),
    .A2(_06123_),
    .B1(_06134_),
    .C1(_06135_),
    .X(_00780_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26679_ (.A(_06124_),
    .X(_06136_));
 sky130_fd_sc_hd__buf_1 _26680_ (.A(_06121_),
    .X(_06137_));
 sky130_fd_sc_hd__a21bo_1 _26681_ (.A1(_06136_),
    .A2(_08265_),
    .B1_N(_06137_),
    .X(_06138_));
 sky130_fd_sc_hd__o211a_1 _26682_ (.A1(net94),
    .A2(_06123_),
    .B1(_06138_),
    .C1(_06135_),
    .X(_00781_));
 sky130_fd_sc_hd__clkbuf_2 _26683_ (.A(_06122_),
    .X(_06139_));
 sky130_fd_sc_hd__a21bo_1 _26684_ (.A1(_06136_),
    .A2(_08266_),
    .B1_N(_06137_),
    .X(_06140_));
 sky130_fd_sc_hd__o211a_1 _26685_ (.A1(net95),
    .A2(_06139_),
    .B1(_06140_),
    .C1(_06135_),
    .X(_00782_));
 sky130_fd_sc_hd__a21bo_1 _26686_ (.A1(_06136_),
    .A2(_08273_),
    .B1_N(_06137_),
    .X(_06141_));
 sky130_fd_sc_hd__o211a_1 _26687_ (.A1(net96),
    .A2(_06139_),
    .B1(_06141_),
    .C1(_06135_),
    .X(_00783_));
 sky130_fd_sc_hd__a21bo_1 _26688_ (.A1(_06136_),
    .A2(_08237_),
    .B1_N(_06137_),
    .X(_06142_));
 sky130_fd_sc_hd__o211a_1 _26689_ (.A1(net97),
    .A2(_06139_),
    .B1(_06142_),
    .C1(_06135_),
    .X(_00784_));
 sky130_fd_sc_hd__a21bo_1 _26690_ (.A1(_06136_),
    .A2(_08252_),
    .B1_N(_06137_),
    .X(_06143_));
 sky130_fd_sc_hd__o211a_1 _26691_ (.A1(net98),
    .A2(_06139_),
    .B1(_06143_),
    .C1(_06135_),
    .X(_00785_));
 sky130_fd_sc_hd__a21bo_1 _26692_ (.A1(_06136_),
    .A2(_08247_),
    .B1_N(_06137_),
    .X(_06144_));
 sky130_fd_sc_hd__clkbuf_2 _26693_ (.A(_06114_),
    .X(_06145_));
 sky130_fd_sc_hd__o211a_1 _26694_ (.A1(net68),
    .A2(_06139_),
    .B1(_06144_),
    .C1(_06145_),
    .X(_00786_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26695_ (.A(_06124_),
    .X(_06146_));
 sky130_fd_sc_hd__buf_1 _26696_ (.A(_06121_),
    .X(_06147_));
 sky130_fd_sc_hd__a21bo_1 _26697_ (.A1(_06146_),
    .A2(_08235_),
    .B1_N(_06147_),
    .X(_06148_));
 sky130_fd_sc_hd__o211a_1 _26698_ (.A1(net69),
    .A2(_06139_),
    .B1(_06148_),
    .C1(_06145_),
    .X(_00787_));
 sky130_fd_sc_hd__clkbuf_2 _26699_ (.A(_06122_),
    .X(_06149_));
 sky130_fd_sc_hd__a21bo_1 _26700_ (.A1(_06146_),
    .A2(_08251_),
    .B1_N(_06147_),
    .X(_06150_));
 sky130_fd_sc_hd__o211a_1 _26701_ (.A1(net70),
    .A2(_06149_),
    .B1(_06150_),
    .C1(_06145_),
    .X(_00788_));
 sky130_fd_sc_hd__a21bo_1 _26702_ (.A1(_06146_),
    .A2(_08260_),
    .B1_N(_06147_),
    .X(_06151_));
 sky130_fd_sc_hd__o211a_1 _26703_ (.A1(net71),
    .A2(_06149_),
    .B1(_06151_),
    .C1(_06145_),
    .X(_00789_));
 sky130_fd_sc_hd__a21bo_1 _26704_ (.A1(_06146_),
    .A2(_08271_),
    .B1_N(_06147_),
    .X(_06152_));
 sky130_fd_sc_hd__o211a_1 _26705_ (.A1(net72),
    .A2(_06149_),
    .B1(_06152_),
    .C1(_06145_),
    .X(_00790_));
 sky130_fd_sc_hd__a21bo_1 _26706_ (.A1(_06146_),
    .A2(_08250_),
    .B1_N(_06147_),
    .X(_06153_));
 sky130_fd_sc_hd__o211a_1 _26707_ (.A1(net73),
    .A2(_06149_),
    .B1(_06153_),
    .C1(_06145_),
    .X(_00791_));
 sky130_fd_sc_hd__a21bo_1 _26708_ (.A1(_06146_),
    .A2(_08257_),
    .B1_N(_06147_),
    .X(_06154_));
 sky130_fd_sc_hd__clkbuf_2 _26709_ (.A(_06114_),
    .X(_06155_));
 sky130_fd_sc_hd__o211a_1 _26710_ (.A1(net74),
    .A2(_06149_),
    .B1(_06154_),
    .C1(_06155_),
    .X(_00792_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26711_ (.A(_06124_),
    .X(_06156_));
 sky130_fd_sc_hd__buf_1 _26712_ (.A(_06120_),
    .X(_06157_));
 sky130_fd_sc_hd__a21bo_1 _26713_ (.A1(_06156_),
    .A2(_08272_),
    .B1_N(_06157_),
    .X(_06158_));
 sky130_fd_sc_hd__o211a_1 _26714_ (.A1(net75),
    .A2(_06149_),
    .B1(_06158_),
    .C1(_06155_),
    .X(_00793_));
 sky130_fd_sc_hd__clkbuf_2 _26715_ (.A(_06122_),
    .X(_06159_));
 sky130_fd_sc_hd__a21bo_1 _26716_ (.A1(_06156_),
    .A2(_08234_),
    .B1_N(_06157_),
    .X(_06160_));
 sky130_fd_sc_hd__o211a_1 _26717_ (.A1(net76),
    .A2(_06159_),
    .B1(_06160_),
    .C1(_06155_),
    .X(_00794_));
 sky130_fd_sc_hd__a21bo_1 _26718_ (.A1(_06156_),
    .A2(_08255_),
    .B1_N(_06157_),
    .X(_06161_));
 sky130_fd_sc_hd__o211a_1 _26719_ (.A1(net77),
    .A2(_06159_),
    .B1(_06161_),
    .C1(_06155_),
    .X(_00795_));
 sky130_fd_sc_hd__a21bo_1 _26720_ (.A1(_06156_),
    .A2(_08244_),
    .B1_N(_06157_),
    .X(_06162_));
 sky130_fd_sc_hd__o211a_1 _26721_ (.A1(net79),
    .A2(_06159_),
    .B1(_06162_),
    .C1(_06155_),
    .X(_00796_));
 sky130_fd_sc_hd__a21bo_1 _26722_ (.A1(_06156_),
    .A2(_08246_),
    .B1_N(_06157_),
    .X(_06163_));
 sky130_fd_sc_hd__o211a_1 _26723_ (.A1(net80),
    .A2(_06159_),
    .B1(_06163_),
    .C1(_06155_),
    .X(_00797_));
 sky130_fd_sc_hd__a21bo_1 _26724_ (.A1(_06156_),
    .A2(_08245_),
    .B1_N(_06157_),
    .X(_06164_));
 sky130_fd_sc_hd__clkbuf_2 _26725_ (.A(_06114_),
    .X(_06165_));
 sky130_fd_sc_hd__o211a_1 _26726_ (.A1(net81),
    .A2(_06159_),
    .B1(_06164_),
    .C1(_06165_),
    .X(_00798_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26727_ (.A(_06124_),
    .X(_06166_));
 sky130_fd_sc_hd__buf_1 _26728_ (.A(_06120_),
    .X(_06167_));
 sky130_fd_sc_hd__a21bo_1 _26729_ (.A1(_06166_),
    .A2(_08249_),
    .B1_N(_06167_),
    .X(_06168_));
 sky130_fd_sc_hd__o211a_1 _26730_ (.A1(net82),
    .A2(_06159_),
    .B1(_06168_),
    .C1(_06165_),
    .X(_00799_));
 sky130_fd_sc_hd__clkbuf_2 _26731_ (.A(_06127_),
    .X(_06169_));
 sky130_fd_sc_hd__a21bo_1 _26732_ (.A1(_06166_),
    .A2(_08262_),
    .B1_N(_06167_),
    .X(_06170_));
 sky130_fd_sc_hd__o211a_1 _26733_ (.A1(net83),
    .A2(_06169_),
    .B1(_06170_),
    .C1(_06165_),
    .X(_00800_));
 sky130_fd_sc_hd__a21bo_1 _26734_ (.A1(_06166_),
    .A2(_08239_),
    .B1_N(_06167_),
    .X(_06171_));
 sky130_fd_sc_hd__o211a_1 _26735_ (.A1(net84),
    .A2(_06169_),
    .B1(_06171_),
    .C1(_06165_),
    .X(_00801_));
 sky130_fd_sc_hd__a21bo_1 _26736_ (.A1(_06166_),
    .A2(_08241_),
    .B1_N(_06167_),
    .X(_06172_));
 sky130_fd_sc_hd__o211a_1 _26737_ (.A1(net85),
    .A2(_06169_),
    .B1(_06172_),
    .C1(_06165_),
    .X(_00802_));
 sky130_fd_sc_hd__a21bo_1 _26738_ (.A1(_06166_),
    .A2(_08261_),
    .B1_N(_06167_),
    .X(_06173_));
 sky130_fd_sc_hd__o211a_1 _26739_ (.A1(net86),
    .A2(_06169_),
    .B1(_06173_),
    .C1(_06165_),
    .X(_00803_));
 sky130_fd_sc_hd__a21bo_1 _26740_ (.A1(_06166_),
    .A2(_08256_),
    .B1_N(_06167_),
    .X(_06174_));
 sky130_fd_sc_hd__buf_2 _26741_ (.A(_06129_),
    .X(_06175_));
 sky130_fd_sc_hd__o211a_1 _26742_ (.A1(net87),
    .A2(_06169_),
    .B1(_06174_),
    .C1(_06175_),
    .X(_00804_));
 sky130_fd_sc_hd__a21bo_1 _26743_ (.A1(_06125_),
    .A2(_08242_),
    .B1_N(_06121_),
    .X(_06176_));
 sky130_fd_sc_hd__o211a_1 _26744_ (.A1(net88),
    .A2(_06169_),
    .B1(_06176_),
    .C1(_06175_),
    .X(_00805_));
 sky130_fd_sc_hd__a21bo_1 _26745_ (.A1(_06125_),
    .A2(_08270_),
    .B1_N(_06121_),
    .X(_06177_));
 sky130_fd_sc_hd__o211a_1 _26746_ (.A1(net90),
    .A2(_06122_),
    .B1(_06177_),
    .C1(_06175_),
    .X(_00806_));
 sky130_fd_sc_hd__a21bo_1 _26747_ (.A1(_06125_),
    .A2(_08258_),
    .B1_N(_06121_),
    .X(_06178_));
 sky130_fd_sc_hd__o211a_1 _26748_ (.A1(net91),
    .A2(_06122_),
    .B1(_06178_),
    .C1(_06175_),
    .X(_00807_));
 sky130_fd_sc_hd__buf_2 _26749_ (.A(_08328_),
    .X(_06179_));
 sky130_fd_sc_hd__clkbuf_4 _26750_ (.A(_06179_),
    .X(_06180_));
 sky130_fd_sc_hd__and2_1 _26751_ (.A(_06180_),
    .B(\cpu_state[0] ),
    .X(_06181_));
 sky130_fd_sc_hd__clkbuf_1 _26752_ (.A(_06181_),
    .X(_00808_));
 sky130_fd_sc_hd__nor2_2 _26753_ (.A(_06117_),
    .B(_08279_),
    .Y(_06182_));
 sky130_fd_sc_hd__and2_1 _26754_ (.A(\count_instr[0] ),
    .B(_06182_),
    .X(_06183_));
 sky130_fd_sc_hd__buf_2 _26755_ (.A(_06179_),
    .X(_06184_));
 sky130_fd_sc_hd__o21ai_1 _26756_ (.A1(\count_instr[0] ),
    .A2(_06182_),
    .B1(_06184_),
    .Y(_06185_));
 sky130_fd_sc_hd__nor2_1 _26757_ (.A(_06183_),
    .B(_06185_),
    .Y(_00809_));
 sky130_fd_sc_hd__and3_1 _26758_ (.A(\count_instr[1] ),
    .B(\count_instr[0] ),
    .C(_06182_),
    .X(_06186_));
 sky130_vsdinv _26759_ (.A(_06186_),
    .Y(_06187_));
 sky130_fd_sc_hd__o211a_1 _26760_ (.A1(\count_instr[1] ),
    .A2(_06183_),
    .B1(_06187_),
    .C1(_06175_),
    .X(_00810_));
 sky130_vsdinv _26761_ (.A(\count_instr[2] ),
    .Y(_06188_));
 sky130_fd_sc_hd__nand2_1 _26762_ (.A(\count_instr[1] ),
    .B(\count_instr[0] ),
    .Y(_06189_));
 sky130_fd_sc_hd__nor4_1 _26763_ (.A(_08145_),
    .B(_06188_),
    .C(_08279_),
    .D(_06189_),
    .Y(_06190_));
 sky130_fd_sc_hd__nor2_1 _26764_ (.A(_08520_),
    .B(_06190_),
    .Y(_06191_));
 sky130_fd_sc_hd__o21a_1 _26765_ (.A1(\count_instr[2] ),
    .A2(_06186_),
    .B1(_06191_),
    .X(_00811_));
 sky130_fd_sc_hd__and2_1 _26766_ (.A(\count_instr[3] ),
    .B(net367),
    .X(_06192_));
 sky130_fd_sc_hd__o21ai_1 _26767_ (.A1(\count_instr[3] ),
    .A2(net367),
    .B1(_06184_),
    .Y(_06193_));
 sky130_fd_sc_hd__nor2_1 _26768_ (.A(_06192_),
    .B(_06193_),
    .Y(_00812_));
 sky130_fd_sc_hd__or2_1 _26769_ (.A(\count_instr[4] ),
    .B(_06192_),
    .X(_06194_));
 sky130_fd_sc_hd__nand2_1 _26770_ (.A(\count_instr[4] ),
    .B(_06192_),
    .Y(_06195_));
 sky130_fd_sc_hd__and3_1 _26771_ (.A(_06129_),
    .B(_06194_),
    .C(_06195_),
    .X(_06196_));
 sky130_fd_sc_hd__clkbuf_1 _26772_ (.A(_06196_),
    .X(_00813_));
 sky130_vsdinv _26773_ (.A(\count_instr[5] ),
    .Y(_06197_));
 sky130_fd_sc_hd__and2_1 _26774_ (.A(\count_instr[5] ),
    .B(\count_instr[4] ),
    .X(_06198_));
 sky130_fd_sc_hd__and3_1 _26775_ (.A(\count_instr[3] ),
    .B(net367),
    .C(_06198_),
    .X(_06199_));
 sky130_fd_sc_hd__buf_2 _26776_ (.A(_08182_),
    .X(_06200_));
 sky130_fd_sc_hd__buf_2 _26777_ (.A(_06200_),
    .X(_06201_));
 sky130_fd_sc_hd__a211oi_1 _26778_ (.A1(_06197_),
    .A2(_06195_),
    .B1(_06199_),
    .C1(_06201_),
    .Y(_00814_));
 sky130_fd_sc_hd__and4_1 _26779_ (.A(\count_instr[6] ),
    .B(\count_instr[3] ),
    .C(net367),
    .D(_06198_),
    .X(_06202_));
 sky130_fd_sc_hd__o21ai_1 _26780_ (.A1(\count_instr[6] ),
    .A2(_06199_),
    .B1(_06184_),
    .Y(_06203_));
 sky130_fd_sc_hd__nor2_1 _26781_ (.A(_06202_),
    .B(_06203_),
    .Y(_00815_));
 sky130_fd_sc_hd__and2_1 _26782_ (.A(\count_instr[7] ),
    .B(_06202_),
    .X(_06204_));
 sky130_fd_sc_hd__clkbuf_2 _26783_ (.A(_08322_),
    .X(_06205_));
 sky130_fd_sc_hd__o21ai_1 _26784_ (.A1(\count_instr[7] ),
    .A2(_06202_),
    .B1(_06205_),
    .Y(_06206_));
 sky130_fd_sc_hd__nor2_1 _26785_ (.A(_06204_),
    .B(_06206_),
    .Y(_00816_));
 sky130_fd_sc_hd__and3_1 _26786_ (.A(\count_instr[8] ),
    .B(\count_instr[7] ),
    .C(_06202_),
    .X(_06207_));
 sky130_fd_sc_hd__o21ai_1 _26787_ (.A1(\count_instr[8] ),
    .A2(_06204_),
    .B1(_06205_),
    .Y(_06208_));
 sky130_fd_sc_hd__nor2_1 _26788_ (.A(_06207_),
    .B(_06208_),
    .Y(_00817_));
 sky130_fd_sc_hd__and4_1 _26789_ (.A(\count_instr[9] ),
    .B(\count_instr[8] ),
    .C(\count_instr[7] ),
    .D(_06202_),
    .X(_06209_));
 sky130_fd_sc_hd__o21ai_1 _26790_ (.A1(\count_instr[9] ),
    .A2(_06207_),
    .B1(_06205_),
    .Y(_06210_));
 sky130_fd_sc_hd__nor2_1 _26791_ (.A(_06209_),
    .B(_06210_),
    .Y(_00818_));
 sky130_fd_sc_hd__a21oi_1 _26792_ (.A1(\count_instr[10] ),
    .A2(_06209_),
    .B1(_06201_),
    .Y(_06211_));
 sky130_fd_sc_hd__o21a_1 _26793_ (.A1(\count_instr[10] ),
    .A2(_06209_),
    .B1(_06211_),
    .X(_00819_));
 sky130_fd_sc_hd__and3_1 _26794_ (.A(\count_instr[11] ),
    .B(\count_instr[10] ),
    .C(_06209_),
    .X(_06212_));
 sky130_fd_sc_hd__a21o_1 _26795_ (.A1(\count_instr[10] ),
    .A2(_06209_),
    .B1(\count_instr[11] ),
    .X(_06213_));
 sky130_fd_sc_hd__and3b_1 _26796_ (.A_N(_06212_),
    .B(_08506_),
    .C(_06213_),
    .X(_06214_));
 sky130_fd_sc_hd__clkbuf_1 _26797_ (.A(_06214_),
    .X(_00820_));
 sky130_fd_sc_hd__and4_1 _26798_ (.A(\count_instr[12] ),
    .B(\count_instr[11] ),
    .C(\count_instr[10] ),
    .D(_06209_),
    .X(_06215_));
 sky130_fd_sc_hd__o21ai_1 _26799_ (.A1(\count_instr[12] ),
    .A2(_06212_),
    .B1(_06205_),
    .Y(_06216_));
 sky130_fd_sc_hd__nor2_1 _26800_ (.A(_06215_),
    .B(_06216_),
    .Y(_00821_));
 sky130_fd_sc_hd__a21oi_1 _26801_ (.A1(\count_instr[13] ),
    .A2(_06215_),
    .B1(_06201_),
    .Y(_06217_));
 sky130_fd_sc_hd__o21a_1 _26802_ (.A1(\count_instr[13] ),
    .A2(_06215_),
    .B1(_06217_),
    .X(_00822_));
 sky130_fd_sc_hd__and3_1 _26803_ (.A(\count_instr[14] ),
    .B(\count_instr[13] ),
    .C(_06215_),
    .X(_06218_));
 sky130_fd_sc_hd__a21o_1 _26804_ (.A1(\count_instr[13] ),
    .A2(_06215_),
    .B1(\count_instr[14] ),
    .X(_06219_));
 sky130_fd_sc_hd__and3b_1 _26805_ (.A_N(_06218_),
    .B(_08506_),
    .C(_06219_),
    .X(_06220_));
 sky130_fd_sc_hd__clkbuf_1 _26806_ (.A(_06220_),
    .X(_00823_));
 sky130_fd_sc_hd__and4_1 _26807_ (.A(\count_instr[15] ),
    .B(\count_instr[14] ),
    .C(\count_instr[13] ),
    .D(_06215_),
    .X(_06221_));
 sky130_fd_sc_hd__o21ai_1 _26808_ (.A1(\count_instr[15] ),
    .A2(_06218_),
    .B1(_06205_),
    .Y(_06222_));
 sky130_fd_sc_hd__nor2_1 _26809_ (.A(_06221_),
    .B(_06222_),
    .Y(_00824_));
 sky130_fd_sc_hd__a21oi_1 _26810_ (.A1(\count_instr[16] ),
    .A2(_06221_),
    .B1(_06201_),
    .Y(_06223_));
 sky130_fd_sc_hd__o21a_1 _26811_ (.A1(\count_instr[16] ),
    .A2(_06221_),
    .B1(_06223_),
    .X(_00825_));
 sky130_fd_sc_hd__and3_1 _26812_ (.A(\count_instr[17] ),
    .B(\count_instr[16] ),
    .C(_06221_),
    .X(_06224_));
 sky130_fd_sc_hd__a21o_1 _26813_ (.A1(\count_instr[16] ),
    .A2(_06221_),
    .B1(\count_instr[17] ),
    .X(_06225_));
 sky130_fd_sc_hd__and3b_1 _26814_ (.A_N(_06224_),
    .B(_08506_),
    .C(_06225_),
    .X(_06226_));
 sky130_fd_sc_hd__clkbuf_1 _26815_ (.A(_06226_),
    .X(_00826_));
 sky130_fd_sc_hd__and4_2 _26816_ (.A(\count_instr[18] ),
    .B(\count_instr[17] ),
    .C(\count_instr[16] ),
    .D(_06221_),
    .X(_06227_));
 sky130_fd_sc_hd__o21ai_1 _26817_ (.A1(\count_instr[18] ),
    .A2(_06224_),
    .B1(_06205_),
    .Y(_06228_));
 sky130_fd_sc_hd__nor2_1 _26818_ (.A(_06227_),
    .B(_06228_),
    .Y(_00827_));
 sky130_fd_sc_hd__buf_2 _26819_ (.A(_06200_),
    .X(_06229_));
 sky130_fd_sc_hd__a21oi_1 _26820_ (.A1(\count_instr[19] ),
    .A2(_06227_),
    .B1(_06229_),
    .Y(_06230_));
 sky130_fd_sc_hd__o21a_1 _26821_ (.A1(\count_instr[19] ),
    .A2(_06227_),
    .B1(_06230_),
    .X(_00828_));
 sky130_fd_sc_hd__and3_1 _26822_ (.A(\count_instr[20] ),
    .B(\count_instr[19] ),
    .C(_06227_),
    .X(_06231_));
 sky130_fd_sc_hd__a21o_1 _26823_ (.A1(\count_instr[19] ),
    .A2(_06227_),
    .B1(\count_instr[20] ),
    .X(_06232_));
 sky130_fd_sc_hd__and3b_1 _26824_ (.A_N(_06231_),
    .B(_08506_),
    .C(_06232_),
    .X(_06233_));
 sky130_fd_sc_hd__clkbuf_1 _26825_ (.A(_06233_),
    .X(_00829_));
 sky130_fd_sc_hd__and4_1 _26826_ (.A(\count_instr[21] ),
    .B(\count_instr[20] ),
    .C(\count_instr[19] ),
    .D(_06227_),
    .X(_06234_));
 sky130_fd_sc_hd__clkbuf_2 _26827_ (.A(_08321_),
    .X(_06235_));
 sky130_fd_sc_hd__clkbuf_2 _26828_ (.A(_06235_),
    .X(_06236_));
 sky130_fd_sc_hd__o21ai_1 _26829_ (.A1(\count_instr[21] ),
    .A2(_06231_),
    .B1(_06236_),
    .Y(_06237_));
 sky130_fd_sc_hd__nor2_1 _26830_ (.A(_06234_),
    .B(_06237_),
    .Y(_00830_));
 sky130_fd_sc_hd__a21oi_1 _26831_ (.A1(\count_instr[22] ),
    .A2(_06234_),
    .B1(_06229_),
    .Y(_06238_));
 sky130_fd_sc_hd__o21a_1 _26832_ (.A1(\count_instr[22] ),
    .A2(_06234_),
    .B1(_06238_),
    .X(_00831_));
 sky130_fd_sc_hd__and3_1 _26833_ (.A(\count_instr[23] ),
    .B(\count_instr[22] ),
    .C(_06234_),
    .X(_06239_));
 sky130_fd_sc_hd__a21o_1 _26834_ (.A1(\count_instr[22] ),
    .A2(_06234_),
    .B1(\count_instr[23] ),
    .X(_06240_));
 sky130_fd_sc_hd__and3b_1 _26835_ (.A_N(_06239_),
    .B(_08506_),
    .C(_06240_),
    .X(_06241_));
 sky130_fd_sc_hd__clkbuf_1 _26836_ (.A(_06241_),
    .X(_00832_));
 sky130_fd_sc_hd__and4_1 _26837_ (.A(\count_instr[24] ),
    .B(\count_instr[23] ),
    .C(\count_instr[22] ),
    .D(_06234_),
    .X(_06242_));
 sky130_fd_sc_hd__o21ai_1 _26838_ (.A1(\count_instr[24] ),
    .A2(_06239_),
    .B1(_06236_),
    .Y(_06243_));
 sky130_fd_sc_hd__nor2_1 _26839_ (.A(_06242_),
    .B(_06243_),
    .Y(_00833_));
 sky130_fd_sc_hd__a21oi_1 _26840_ (.A1(\count_instr[25] ),
    .A2(_06242_),
    .B1(_06229_),
    .Y(_06244_));
 sky130_fd_sc_hd__o21a_1 _26841_ (.A1(\count_instr[25] ),
    .A2(_06242_),
    .B1(_06244_),
    .X(_00834_));
 sky130_fd_sc_hd__and3_1 _26842_ (.A(\count_instr[26] ),
    .B(\count_instr[25] ),
    .C(_06242_),
    .X(_06245_));
 sky130_fd_sc_hd__clkbuf_2 _26843_ (.A(_06179_),
    .X(_06246_));
 sky130_fd_sc_hd__a21o_1 _26844_ (.A1(\count_instr[25] ),
    .A2(_06242_),
    .B1(\count_instr[26] ),
    .X(_06247_));
 sky130_fd_sc_hd__and3b_1 _26845_ (.A_N(_06245_),
    .B(_06246_),
    .C(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__clkbuf_1 _26846_ (.A(_06248_),
    .X(_00835_));
 sky130_fd_sc_hd__and4_1 _26847_ (.A(\count_instr[27] ),
    .B(\count_instr[26] ),
    .C(\count_instr[25] ),
    .D(_06242_),
    .X(_06249_));
 sky130_fd_sc_hd__o21ai_1 _26848_ (.A1(\count_instr[27] ),
    .A2(_06245_),
    .B1(_06236_),
    .Y(_06250_));
 sky130_fd_sc_hd__nor2_1 _26849_ (.A(_06249_),
    .B(_06250_),
    .Y(_00836_));
 sky130_fd_sc_hd__a21oi_1 _26850_ (.A1(\count_instr[28] ),
    .A2(_06249_),
    .B1(_06229_),
    .Y(_06251_));
 sky130_fd_sc_hd__o21a_1 _26851_ (.A1(\count_instr[28] ),
    .A2(_06249_),
    .B1(_06251_),
    .X(_00837_));
 sky130_fd_sc_hd__and3_1 _26852_ (.A(\count_instr[29] ),
    .B(\count_instr[28] ),
    .C(_06249_),
    .X(_06252_));
 sky130_fd_sc_hd__a21o_1 _26853_ (.A1(\count_instr[28] ),
    .A2(_06249_),
    .B1(\count_instr[29] ),
    .X(_06253_));
 sky130_fd_sc_hd__and3b_1 _26854_ (.A_N(_06252_),
    .B(_06246_),
    .C(_06253_),
    .X(_06254_));
 sky130_fd_sc_hd__clkbuf_1 _26855_ (.A(_06254_),
    .X(_00838_));
 sky130_fd_sc_hd__and4_2 _26856_ (.A(\count_instr[30] ),
    .B(\count_instr[29] ),
    .C(\count_instr[28] ),
    .D(_06249_),
    .X(_06255_));
 sky130_fd_sc_hd__o21ai_1 _26857_ (.A1(\count_instr[30] ),
    .A2(_06252_),
    .B1(_06236_),
    .Y(_06256_));
 sky130_fd_sc_hd__nor2_1 _26858_ (.A(_06255_),
    .B(_06256_),
    .Y(_00839_));
 sky130_fd_sc_hd__a21oi_1 _26859_ (.A1(\count_instr[31] ),
    .A2(_06255_),
    .B1(_06229_),
    .Y(_06257_));
 sky130_fd_sc_hd__o21a_1 _26860_ (.A1(\count_instr[31] ),
    .A2(_06255_),
    .B1(_06257_),
    .X(_00840_));
 sky130_fd_sc_hd__and3_1 _26861_ (.A(\count_instr[32] ),
    .B(\count_instr[31] ),
    .C(_06255_),
    .X(_06258_));
 sky130_fd_sc_hd__a21o_1 _26862_ (.A1(\count_instr[31] ),
    .A2(_06255_),
    .B1(\count_instr[32] ),
    .X(_06259_));
 sky130_fd_sc_hd__and3b_1 _26863_ (.A_N(_06258_),
    .B(_06246_),
    .C(_06259_),
    .X(_06260_));
 sky130_fd_sc_hd__clkbuf_1 _26864_ (.A(_06260_),
    .X(_00841_));
 sky130_fd_sc_hd__or2_1 _26865_ (.A(\count_instr[33] ),
    .B(_06258_),
    .X(_06261_));
 sky130_fd_sc_hd__nand2_1 _26866_ (.A(\count_instr[33] ),
    .B(_06258_),
    .Y(_06262_));
 sky130_fd_sc_hd__and3_1 _26867_ (.A(_06129_),
    .B(_06261_),
    .C(_06262_),
    .X(_06263_));
 sky130_fd_sc_hd__clkbuf_1 _26868_ (.A(_06263_),
    .X(_00842_));
 sky130_vsdinv _26869_ (.A(\count_instr[34] ),
    .Y(_06264_));
 sky130_fd_sc_hd__and2_1 _26870_ (.A(\count_instr[34] ),
    .B(\count_instr[33] ),
    .X(_06265_));
 sky130_fd_sc_hd__and4_1 _26871_ (.A(\count_instr[32] ),
    .B(\count_instr[31] ),
    .C(_06255_),
    .D(_06265_),
    .X(_06266_));
 sky130_fd_sc_hd__a211oi_1 _26872_ (.A1(_06264_),
    .A2(_06262_),
    .B1(_06266_),
    .C1(_06201_),
    .Y(_00843_));
 sky130_fd_sc_hd__and2_1 _26873_ (.A(\count_instr[35] ),
    .B(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__o21ai_1 _26874_ (.A1(\count_instr[35] ),
    .A2(_06266_),
    .B1(_06236_),
    .Y(_06268_));
 sky130_fd_sc_hd__nor2_1 _26875_ (.A(_06267_),
    .B(_06268_),
    .Y(_00844_));
 sky130_fd_sc_hd__and3_1 _26876_ (.A(\count_instr[36] ),
    .B(\count_instr[35] ),
    .C(_06266_),
    .X(_06269_));
 sky130_fd_sc_hd__o21ai_1 _26877_ (.A1(\count_instr[36] ),
    .A2(_06267_),
    .B1(_06236_),
    .Y(_06270_));
 sky130_fd_sc_hd__nor2_1 _26878_ (.A(_06269_),
    .B(_06270_),
    .Y(_00845_));
 sky130_fd_sc_hd__and4_1 _26879_ (.A(\count_instr[37] ),
    .B(\count_instr[36] ),
    .C(\count_instr[35] ),
    .D(_06266_),
    .X(_06271_));
 sky130_fd_sc_hd__clkbuf_2 _26880_ (.A(_06235_),
    .X(_06272_));
 sky130_fd_sc_hd__o21ai_1 _26881_ (.A1(\count_instr[37] ),
    .A2(_06269_),
    .B1(_06272_),
    .Y(_06273_));
 sky130_fd_sc_hd__nor2_1 _26882_ (.A(_06271_),
    .B(_06273_),
    .Y(_00846_));
 sky130_fd_sc_hd__and2_1 _26883_ (.A(\count_instr[38] ),
    .B(_06271_),
    .X(_06274_));
 sky130_fd_sc_hd__o21ai_1 _26884_ (.A1(\count_instr[38] ),
    .A2(_06271_),
    .B1(_06272_),
    .Y(_06275_));
 sky130_fd_sc_hd__nor2_1 _26885_ (.A(_06274_),
    .B(_06275_),
    .Y(_00847_));
 sky130_fd_sc_hd__and3_1 _26886_ (.A(\count_instr[39] ),
    .B(\count_instr[38] ),
    .C(_06271_),
    .X(_06276_));
 sky130_fd_sc_hd__o21ai_1 _26887_ (.A1(\count_instr[39] ),
    .A2(_06274_),
    .B1(_06272_),
    .Y(_06277_));
 sky130_fd_sc_hd__nor2_1 _26888_ (.A(_06276_),
    .B(_06277_),
    .Y(_00848_));
 sky130_fd_sc_hd__and4_1 _26889_ (.A(\count_instr[40] ),
    .B(\count_instr[39] ),
    .C(\count_instr[38] ),
    .D(_06271_),
    .X(_06278_));
 sky130_fd_sc_hd__o21ai_1 _26890_ (.A1(\count_instr[40] ),
    .A2(_06276_),
    .B1(_06272_),
    .Y(_06279_));
 sky130_fd_sc_hd__nor2_1 _26891_ (.A(_06278_),
    .B(_06279_),
    .Y(_00849_));
 sky130_fd_sc_hd__a21oi_1 _26892_ (.A1(\count_instr[41] ),
    .A2(_06278_),
    .B1(_06229_),
    .Y(_06280_));
 sky130_fd_sc_hd__o21a_1 _26893_ (.A1(\count_instr[41] ),
    .A2(_06278_),
    .B1(_06280_),
    .X(_00850_));
 sky130_fd_sc_hd__and3_1 _26894_ (.A(\count_instr[42] ),
    .B(\count_instr[41] ),
    .C(_06278_),
    .X(_06281_));
 sky130_fd_sc_hd__a21o_1 _26895_ (.A1(\count_instr[41] ),
    .A2(_06278_),
    .B1(\count_instr[42] ),
    .X(_06282_));
 sky130_fd_sc_hd__and3b_1 _26896_ (.A_N(_06281_),
    .B(_06246_),
    .C(_06282_),
    .X(_06283_));
 sky130_fd_sc_hd__clkbuf_1 _26897_ (.A(_06283_),
    .X(_00851_));
 sky130_fd_sc_hd__and4_2 _26898_ (.A(\count_instr[43] ),
    .B(\count_instr[42] ),
    .C(\count_instr[41] ),
    .D(_06278_),
    .X(_06284_));
 sky130_fd_sc_hd__o21ai_1 _26899_ (.A1(\count_instr[43] ),
    .A2(_06281_),
    .B1(_06272_),
    .Y(_06285_));
 sky130_fd_sc_hd__nor2_1 _26900_ (.A(_06284_),
    .B(_06285_),
    .Y(_00852_));
 sky130_fd_sc_hd__buf_2 _26901_ (.A(_06200_),
    .X(_06286_));
 sky130_fd_sc_hd__a21oi_1 _26902_ (.A1(\count_instr[44] ),
    .A2(_06284_),
    .B1(_06286_),
    .Y(_06287_));
 sky130_fd_sc_hd__o21a_1 _26903_ (.A1(\count_instr[44] ),
    .A2(_06284_),
    .B1(_06287_),
    .X(_00853_));
 sky130_fd_sc_hd__and3_1 _26904_ (.A(\count_instr[45] ),
    .B(\count_instr[44] ),
    .C(_06284_),
    .X(_06288_));
 sky130_fd_sc_hd__a21o_1 _26905_ (.A1(\count_instr[44] ),
    .A2(_06284_),
    .B1(\count_instr[45] ),
    .X(_06289_));
 sky130_fd_sc_hd__and3b_1 _26906_ (.A_N(_06288_),
    .B(_06246_),
    .C(_06289_),
    .X(_06290_));
 sky130_fd_sc_hd__clkbuf_1 _26907_ (.A(_06290_),
    .X(_00854_));
 sky130_fd_sc_hd__and4_2 _26908_ (.A(\count_instr[46] ),
    .B(\count_instr[45] ),
    .C(\count_instr[44] ),
    .D(_06284_),
    .X(_06291_));
 sky130_fd_sc_hd__o21ai_1 _26909_ (.A1(\count_instr[46] ),
    .A2(_06288_),
    .B1(_06272_),
    .Y(_06292_));
 sky130_fd_sc_hd__nor2_1 _26910_ (.A(_06291_),
    .B(_06292_),
    .Y(_00855_));
 sky130_fd_sc_hd__a21oi_1 _26911_ (.A1(\count_instr[47] ),
    .A2(_06291_),
    .B1(_06286_),
    .Y(_06293_));
 sky130_fd_sc_hd__o21a_1 _26912_ (.A1(\count_instr[47] ),
    .A2(_06291_),
    .B1(_06293_),
    .X(_00856_));
 sky130_fd_sc_hd__and3_1 _26913_ (.A(\count_instr[48] ),
    .B(\count_instr[47] ),
    .C(_06291_),
    .X(_06294_));
 sky130_fd_sc_hd__a21o_1 _26914_ (.A1(\count_instr[47] ),
    .A2(_06291_),
    .B1(\count_instr[48] ),
    .X(_06295_));
 sky130_fd_sc_hd__and3b_1 _26915_ (.A_N(_06294_),
    .B(_06246_),
    .C(_06295_),
    .X(_06296_));
 sky130_fd_sc_hd__clkbuf_1 _26916_ (.A(_06296_),
    .X(_00857_));
 sky130_fd_sc_hd__and4_2 _26917_ (.A(\count_instr[49] ),
    .B(\count_instr[48] ),
    .C(\count_instr[47] ),
    .D(_06291_),
    .X(_06297_));
 sky130_fd_sc_hd__clkbuf_2 _26918_ (.A(_06235_),
    .X(_06298_));
 sky130_fd_sc_hd__o21ai_1 _26919_ (.A1(\count_instr[49] ),
    .A2(_06294_),
    .B1(_06298_),
    .Y(_06299_));
 sky130_fd_sc_hd__nor2_1 _26920_ (.A(_06297_),
    .B(_06299_),
    .Y(_00858_));
 sky130_fd_sc_hd__a21oi_1 _26921_ (.A1(\count_instr[50] ),
    .A2(_06297_),
    .B1(_06286_),
    .Y(_06300_));
 sky130_fd_sc_hd__o21a_1 _26922_ (.A1(\count_instr[50] ),
    .A2(_06297_),
    .B1(_06300_),
    .X(_00859_));
 sky130_fd_sc_hd__and3_1 _26923_ (.A(\count_instr[51] ),
    .B(\count_instr[50] ),
    .C(_06297_),
    .X(_06301_));
 sky130_fd_sc_hd__buf_2 _26924_ (.A(_06179_),
    .X(_06302_));
 sky130_fd_sc_hd__a21o_1 _26925_ (.A1(\count_instr[50] ),
    .A2(_06297_),
    .B1(\count_instr[51] ),
    .X(_06303_));
 sky130_fd_sc_hd__and3b_1 _26926_ (.A_N(_06301_),
    .B(_06302_),
    .C(_06303_),
    .X(_06304_));
 sky130_fd_sc_hd__clkbuf_1 _26927_ (.A(_06304_),
    .X(_00860_));
 sky130_fd_sc_hd__and4_1 _26928_ (.A(\count_instr[52] ),
    .B(\count_instr[51] ),
    .C(\count_instr[50] ),
    .D(_06297_),
    .X(_06305_));
 sky130_fd_sc_hd__o21ai_1 _26929_ (.A1(\count_instr[52] ),
    .A2(_06301_),
    .B1(_06298_),
    .Y(_06306_));
 sky130_fd_sc_hd__nor2_1 _26930_ (.A(_06305_),
    .B(_06306_),
    .Y(_00861_));
 sky130_fd_sc_hd__a21oi_1 _26931_ (.A1(\count_instr[53] ),
    .A2(_06305_),
    .B1(_06286_),
    .Y(_06307_));
 sky130_fd_sc_hd__o21a_1 _26932_ (.A1(\count_instr[53] ),
    .A2(_06305_),
    .B1(_06307_),
    .X(_00862_));
 sky130_fd_sc_hd__and3_1 _26933_ (.A(\count_instr[54] ),
    .B(\count_instr[53] ),
    .C(_06305_),
    .X(_06308_));
 sky130_fd_sc_hd__a21o_1 _26934_ (.A1(\count_instr[53] ),
    .A2(_06305_),
    .B1(\count_instr[54] ),
    .X(_06309_));
 sky130_fd_sc_hd__and3b_1 _26935_ (.A_N(_06308_),
    .B(_06302_),
    .C(_06309_),
    .X(_06310_));
 sky130_fd_sc_hd__clkbuf_1 _26936_ (.A(_06310_),
    .X(_00863_));
 sky130_fd_sc_hd__and4_1 _26937_ (.A(\count_instr[55] ),
    .B(\count_instr[54] ),
    .C(\count_instr[53] ),
    .D(_06305_),
    .X(_06311_));
 sky130_fd_sc_hd__o21ai_1 _26938_ (.A1(\count_instr[55] ),
    .A2(_06308_),
    .B1(_06298_),
    .Y(_06312_));
 sky130_fd_sc_hd__nor2_1 _26939_ (.A(_06311_),
    .B(_06312_),
    .Y(_00864_));
 sky130_fd_sc_hd__and2_1 _26940_ (.A(\count_instr[56] ),
    .B(_06311_),
    .X(_06313_));
 sky130_fd_sc_hd__o21ai_1 _26941_ (.A1(\count_instr[56] ),
    .A2(_06311_),
    .B1(_06298_),
    .Y(_06314_));
 sky130_fd_sc_hd__nor2_1 _26942_ (.A(_06313_),
    .B(_06314_),
    .Y(_00865_));
 sky130_fd_sc_hd__and3_1 _26943_ (.A(\count_instr[57] ),
    .B(\count_instr[56] ),
    .C(_06311_),
    .X(_06315_));
 sky130_fd_sc_hd__o21ai_1 _26944_ (.A1(\count_instr[57] ),
    .A2(_06313_),
    .B1(_06298_),
    .Y(_06316_));
 sky130_fd_sc_hd__nor2_1 _26945_ (.A(_06315_),
    .B(_06316_),
    .Y(_00866_));
 sky130_fd_sc_hd__and2_1 _26946_ (.A(\count_instr[58] ),
    .B(_06315_),
    .X(_06317_));
 sky130_fd_sc_hd__o21ai_1 _26947_ (.A1(\count_instr[58] ),
    .A2(_06315_),
    .B1(_06298_),
    .Y(_06318_));
 sky130_fd_sc_hd__nor2_1 _26948_ (.A(_06317_),
    .B(_06318_),
    .Y(_00867_));
 sky130_fd_sc_hd__a21oi_1 _26949_ (.A1(\count_instr[59] ),
    .A2(_06317_),
    .B1(_06286_),
    .Y(_06319_));
 sky130_fd_sc_hd__o21a_1 _26950_ (.A1(\count_instr[59] ),
    .A2(_06317_),
    .B1(_06319_),
    .X(_00868_));
 sky130_fd_sc_hd__and3_1 _26951_ (.A(\count_instr[60] ),
    .B(\count_instr[59] ),
    .C(_06317_),
    .X(_06320_));
 sky130_fd_sc_hd__a31o_1 _26952_ (.A1(\count_instr[59] ),
    .A2(\count_instr[58] ),
    .A3(_06315_),
    .B1(\count_instr[60] ),
    .X(_06321_));
 sky130_fd_sc_hd__and3b_1 _26953_ (.A_N(_06320_),
    .B(_06302_),
    .C(_06321_),
    .X(_06322_));
 sky130_fd_sc_hd__clkbuf_1 _26954_ (.A(_06322_),
    .X(_00869_));
 sky130_fd_sc_hd__and2_1 _26955_ (.A(\count_instr[61] ),
    .B(_06320_),
    .X(_06323_));
 sky130_fd_sc_hd__buf_2 _26956_ (.A(_06235_),
    .X(_06324_));
 sky130_fd_sc_hd__o21ai_1 _26957_ (.A1(\count_instr[61] ),
    .A2(_06320_),
    .B1(_06324_),
    .Y(_06325_));
 sky130_fd_sc_hd__nor2_1 _26958_ (.A(_06323_),
    .B(_06325_),
    .Y(_00870_));
 sky130_fd_sc_hd__and3_1 _26959_ (.A(\count_instr[62] ),
    .B(\count_instr[61] ),
    .C(_06320_),
    .X(_06326_));
 sky130_fd_sc_hd__o21ai_1 _26960_ (.A1(\count_instr[62] ),
    .A2(_06323_),
    .B1(_06324_),
    .Y(_06327_));
 sky130_fd_sc_hd__nor2_1 _26961_ (.A(_06326_),
    .B(_06327_),
    .Y(_00871_));
 sky130_fd_sc_hd__clkbuf_2 _26962_ (.A(_06179_),
    .X(_06328_));
 sky130_fd_sc_hd__o21ai_1 _26963_ (.A1(\count_instr[63] ),
    .A2(_06326_),
    .B1(_06328_),
    .Y(_06329_));
 sky130_fd_sc_hd__a21oi_1 _26964_ (.A1(\count_instr[63] ),
    .A2(_06326_),
    .B1(_06329_),
    .Y(_00872_));
 sky130_fd_sc_hd__nor2_1 _26965_ (.A(_08232_),
    .B(_08182_),
    .Y(_06330_));
 sky130_fd_sc_hd__buf_2 _26966_ (.A(_06330_),
    .X(_06331_));
 sky130_fd_sc_hd__clkbuf_2 _26967_ (.A(_06331_),
    .X(_06332_));
 sky130_fd_sc_hd__clkbuf_2 _26968_ (.A(_08176_),
    .X(_06333_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26969_ (.A(_06333_),
    .X(_06334_));
 sky130_fd_sc_hd__or2b_2 _26970_ (.A(latched_branch),
    .B_N(\irq_state[0] ),
    .X(_06335_));
 sky130_fd_sc_hd__and2_2 _26971_ (.A(_10313_),
    .B(_06335_),
    .X(_06336_));
 sky130_fd_sc_hd__a22o_2 _26972_ (.A1(_10324_),
    .A2(_05000_),
    .B1(_06336_),
    .B2(\reg_next_pc[1] ),
    .X(_06337_));
 sky130_fd_sc_hd__a22o_1 _26973_ (.A1(_08184_),
    .A2(_06332_),
    .B1(_06334_),
    .B2(_06337_),
    .X(_00873_));
 sky130_fd_sc_hd__o211a_1 _26974_ (.A1(_10312_),
    .A2(_05010_),
    .B1(_06335_),
    .C1(_10318_),
    .X(_06338_));
 sky130_fd_sc_hd__clkbuf_2 _26975_ (.A(_06338_),
    .X(_06339_));
 sky130_fd_sc_hd__a22o_1 _26976_ (.A1(_05008_),
    .A2(_06332_),
    .B1(_06334_),
    .B2(_06339_),
    .X(_00874_));
 sky130_fd_sc_hd__and2_1 _26977_ (.A(_10323_),
    .B(_05018_),
    .X(_06340_));
 sky130_fd_sc_hd__a31o_1 _26978_ (.A1(\reg_next_pc[3] ),
    .A2(_10313_),
    .A3(_06335_),
    .B1(_06340_),
    .X(_06341_));
 sky130_fd_sc_hd__clkbuf_2 _26979_ (.A(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__a22o_1 _26980_ (.A1(_08874_),
    .A2(_06332_),
    .B1(_06334_),
    .B2(_06342_),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _26981_ (.A0(\reg_next_pc[4] ),
    .A1(_05026_),
    .S(_10323_),
    .X(_06343_));
 sky130_fd_sc_hd__or2_1 _26982_ (.A(\irq_state[0] ),
    .B(_06343_),
    .X(_06344_));
 sky130_fd_sc_hd__buf_2 _26983_ (.A(_06344_),
    .X(_06345_));
 sky130_fd_sc_hd__a22o_1 _26984_ (.A1(\reg_pc[4] ),
    .A2(_06332_),
    .B1(_06334_),
    .B2(_06345_),
    .X(_00876_));
 sky130_fd_sc_hd__buf_2 _26985_ (.A(_06330_),
    .X(_06346_));
 sky130_fd_sc_hd__clkbuf_2 _26986_ (.A(_06346_),
    .X(_06347_));
 sky130_fd_sc_hd__a22o_1 _26987_ (.A1(_10324_),
    .A2(_05034_),
    .B1(_06336_),
    .B2(\reg_next_pc[5] ),
    .X(_06348_));
 sky130_fd_sc_hd__clkbuf_2 _26988_ (.A(_06348_),
    .X(_06349_));
 sky130_fd_sc_hd__a22o_1 _26989_ (.A1(\reg_pc[5] ),
    .A2(_06347_),
    .B1(_06334_),
    .B2(_06349_),
    .X(_00877_));
 sky130_fd_sc_hd__and2_1 _26990_ (.A(_10324_),
    .B(_05043_),
    .X(_06350_));
 sky130_fd_sc_hd__a31o_1 _26991_ (.A1(\reg_next_pc[6] ),
    .A2(_10313_),
    .A3(_06335_),
    .B1(_06350_),
    .X(_06351_));
 sky130_fd_sc_hd__clkbuf_2 _26992_ (.A(_06351_),
    .X(_06352_));
 sky130_fd_sc_hd__a22o_1 _26993_ (.A1(_08997_),
    .A2(_06347_),
    .B1(_06334_),
    .B2(_06352_),
    .X(_00878_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26994_ (.A(_06333_),
    .X(_06353_));
 sky130_fd_sc_hd__a22o_1 _26995_ (.A1(_10324_),
    .A2(_05053_),
    .B1(_06336_),
    .B2(\reg_next_pc[7] ),
    .X(_06354_));
 sky130_fd_sc_hd__clkbuf_2 _26996_ (.A(_06354_),
    .X(_06355_));
 sky130_fd_sc_hd__a22o_1 _26997_ (.A1(\reg_pc[7] ),
    .A2(_06347_),
    .B1(_06353_),
    .B2(_06355_),
    .X(_00879_));
 sky130_fd_sc_hd__and3_1 _26998_ (.A(\reg_next_pc[8] ),
    .B(_10313_),
    .C(_06335_),
    .X(_06356_));
 sky130_fd_sc_hd__a21o_1 _26999_ (.A1(_10324_),
    .A2(_05062_),
    .B1(_06356_),
    .X(_06357_));
 sky130_fd_sc_hd__clkbuf_2 _27000_ (.A(_06357_),
    .X(_06358_));
 sky130_fd_sc_hd__a22o_1 _27001_ (.A1(\reg_pc[8] ),
    .A2(_06347_),
    .B1(_06353_),
    .B2(_06358_),
    .X(_00880_));
 sky130_fd_sc_hd__a22o_1 _27002_ (.A1(_10325_),
    .A2(_05072_),
    .B1(_06336_),
    .B2(\reg_next_pc[9] ),
    .X(_06359_));
 sky130_fd_sc_hd__clkbuf_2 _27003_ (.A(_06359_),
    .X(_06360_));
 sky130_fd_sc_hd__a22o_1 _27004_ (.A1(_09170_),
    .A2(_06347_),
    .B1(_06353_),
    .B2(_06360_),
    .X(_00881_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27005_ (.A(_06335_),
    .X(_06361_));
 sky130_fd_sc_hd__o21a_2 _27006_ (.A1(_10316_),
    .A2(_04971_),
    .B1(_10317_),
    .X(_06362_));
 sky130_fd_sc_hd__o22a_1 _27007_ (.A1(_10313_),
    .A2(_05078_),
    .B1(_06362_),
    .B2(\reg_next_pc[10] ),
    .X(_06363_));
 sky130_fd_sc_hd__and2_1 _27008_ (.A(_06361_),
    .B(_06363_),
    .X(_06364_));
 sky130_fd_sc_hd__clkbuf_2 _27009_ (.A(_06364_),
    .X(_06365_));
 sky130_fd_sc_hd__a22o_1 _27010_ (.A1(_09218_),
    .A2(_06347_),
    .B1(_06353_),
    .B2(_06365_),
    .X(_00882_));
 sky130_fd_sc_hd__clkbuf_2 _27011_ (.A(_06346_),
    .X(_06366_));
 sky130_fd_sc_hd__a22o_1 _27012_ (.A1(_10325_),
    .A2(_05087_),
    .B1(_06336_),
    .B2(\reg_next_pc[11] ),
    .X(_06367_));
 sky130_fd_sc_hd__clkbuf_2 _27013_ (.A(_06367_),
    .X(_06368_));
 sky130_fd_sc_hd__a22o_1 _27014_ (.A1(_09295_),
    .A2(_06366_),
    .B1(_06353_),
    .B2(_06368_),
    .X(_00883_));
 sky130_fd_sc_hd__o22a_1 _27015_ (.A1(_10314_),
    .A2(_05098_),
    .B1(_06362_),
    .B2(\reg_next_pc[12] ),
    .X(_06369_));
 sky130_fd_sc_hd__and2_1 _27016_ (.A(_06361_),
    .B(_06369_),
    .X(_06370_));
 sky130_fd_sc_hd__clkbuf_2 _27017_ (.A(_06370_),
    .X(_06371_));
 sky130_fd_sc_hd__a22o_1 _27018_ (.A1(_09347_),
    .A2(_06366_),
    .B1(_06353_),
    .B2(_06371_),
    .X(_00884_));
 sky130_fd_sc_hd__clkbuf_2 _27019_ (.A(_06333_),
    .X(_06372_));
 sky130_fd_sc_hd__clkbuf_2 _27020_ (.A(_06336_),
    .X(_06373_));
 sky130_fd_sc_hd__a22o_1 _27021_ (.A1(_10325_),
    .A2(_05106_),
    .B1(_06373_),
    .B2(\reg_next_pc[13] ),
    .X(_06374_));
 sky130_fd_sc_hd__clkbuf_2 _27022_ (.A(_06374_),
    .X(_06375_));
 sky130_fd_sc_hd__a22o_1 _27023_ (.A1(\reg_pc[13] ),
    .A2(_06366_),
    .B1(_06372_),
    .B2(_06375_),
    .X(_00885_));
 sky130_fd_sc_hd__o22a_1 _27024_ (.A1(_10314_),
    .A2(_05115_),
    .B1(_06362_),
    .B2(\reg_next_pc[14] ),
    .X(_06376_));
 sky130_fd_sc_hd__and2_1 _27025_ (.A(_06361_),
    .B(_06376_),
    .X(_06377_));
 sky130_fd_sc_hd__clkbuf_2 _27026_ (.A(_06377_),
    .X(_06378_));
 sky130_fd_sc_hd__a22o_1 _27027_ (.A1(_09386_),
    .A2(_06366_),
    .B1(_06372_),
    .B2(_06378_),
    .X(_00886_));
 sky130_fd_sc_hd__a22o_1 _27028_ (.A1(_10325_),
    .A2(_05123_),
    .B1(_06373_),
    .B2(\reg_next_pc[15] ),
    .X(_06379_));
 sky130_fd_sc_hd__clkbuf_2 _27029_ (.A(_06379_),
    .X(_06380_));
 sky130_fd_sc_hd__a22o_1 _27030_ (.A1(\reg_pc[15] ),
    .A2(_06366_),
    .B1(_06372_),
    .B2(_06380_),
    .X(_00887_));
 sky130_fd_sc_hd__o22a_1 _27031_ (.A1(_10314_),
    .A2(_05131_),
    .B1(_06362_),
    .B2(\reg_next_pc[16] ),
    .X(_06381_));
 sky130_fd_sc_hd__and2_1 _27032_ (.A(_06361_),
    .B(_06381_),
    .X(_06382_));
 sky130_fd_sc_hd__clkbuf_2 _27033_ (.A(_06382_),
    .X(_06383_));
 sky130_fd_sc_hd__a22o_1 _27034_ (.A1(_09468_),
    .A2(_06366_),
    .B1(_06372_),
    .B2(_06383_),
    .X(_00888_));
 sky130_fd_sc_hd__clkbuf_2 _27035_ (.A(_06346_),
    .X(_06384_));
 sky130_fd_sc_hd__a22o_1 _27036_ (.A1(_10325_),
    .A2(_05140_),
    .B1(_06373_),
    .B2(\reg_next_pc[17] ),
    .X(_06385_));
 sky130_fd_sc_hd__clkbuf_2 _27037_ (.A(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__a22o_1 _27038_ (.A1(\reg_pc[17] ),
    .A2(_06384_),
    .B1(_06372_),
    .B2(_06386_),
    .X(_00889_));
 sky130_fd_sc_hd__o22a_1 _27039_ (.A1(_10314_),
    .A2(_05148_),
    .B1(_06362_),
    .B2(\reg_next_pc[18] ),
    .X(_06387_));
 sky130_fd_sc_hd__and2_1 _27040_ (.A(_06361_),
    .B(_06387_),
    .X(_06388_));
 sky130_fd_sc_hd__clkbuf_2 _27041_ (.A(_06388_),
    .X(_06389_));
 sky130_fd_sc_hd__a22o_1 _27042_ (.A1(_05150_),
    .A2(_06384_),
    .B1(_06372_),
    .B2(_06389_),
    .X(_00890_));
 sky130_fd_sc_hd__buf_2 _27043_ (.A(_08176_),
    .X(_06390_));
 sky130_fd_sc_hd__clkbuf_2 _27044_ (.A(_06390_),
    .X(_06391_));
 sky130_fd_sc_hd__a22o_1 _27045_ (.A1(_10326_),
    .A2(_05158_),
    .B1(_06373_),
    .B2(\reg_next_pc[19] ),
    .X(_06392_));
 sky130_fd_sc_hd__clkbuf_2 _27046_ (.A(_06392_),
    .X(_06393_));
 sky130_fd_sc_hd__a22o_1 _27047_ (.A1(\reg_pc[19] ),
    .A2(_06384_),
    .B1(_06391_),
    .B2(_06393_),
    .X(_00891_));
 sky130_fd_sc_hd__clkbuf_2 _27048_ (.A(_06361_),
    .X(_06394_));
 sky130_fd_sc_hd__clkbuf_2 _27049_ (.A(_06362_),
    .X(_06395_));
 sky130_fd_sc_hd__o22a_1 _27050_ (.A1(_10314_),
    .A2(_05167_),
    .B1(_06395_),
    .B2(\reg_next_pc[20] ),
    .X(_06396_));
 sky130_fd_sc_hd__and2_1 _27051_ (.A(_06394_),
    .B(_06396_),
    .X(_06397_));
 sky130_fd_sc_hd__clkbuf_2 _27052_ (.A(_06397_),
    .X(_06398_));
 sky130_fd_sc_hd__a22o_1 _27053_ (.A1(_09634_),
    .A2(_06384_),
    .B1(_06391_),
    .B2(_06398_),
    .X(_00892_));
 sky130_fd_sc_hd__a22o_2 _27054_ (.A1(_10326_),
    .A2(_05175_),
    .B1(_06373_),
    .B2(\reg_next_pc[21] ),
    .X(_06399_));
 sky130_fd_sc_hd__clkbuf_2 _27055_ (.A(_06399_),
    .X(_06400_));
 sky130_fd_sc_hd__a22o_1 _27056_ (.A1(\reg_pc[21] ),
    .A2(_06384_),
    .B1(_06391_),
    .B2(_06400_),
    .X(_00893_));
 sky130_fd_sc_hd__o22a_1 _27057_ (.A1(_10315_),
    .A2(_05184_),
    .B1(_06395_),
    .B2(\reg_next_pc[22] ),
    .X(_06401_));
 sky130_fd_sc_hd__and2_1 _27058_ (.A(_06394_),
    .B(_06401_),
    .X(_06402_));
 sky130_fd_sc_hd__clkbuf_2 _27059_ (.A(_06402_),
    .X(_06403_));
 sky130_fd_sc_hd__a22o_1 _27060_ (.A1(_09712_),
    .A2(_06384_),
    .B1(_06391_),
    .B2(_06403_),
    .X(_00894_));
 sky130_fd_sc_hd__clkbuf_2 _27061_ (.A(_06331_),
    .X(_06404_));
 sky130_fd_sc_hd__buf_2 _27062_ (.A(_06373_),
    .X(_06405_));
 sky130_fd_sc_hd__a22o_1 _27063_ (.A1(_10326_),
    .A2(_05193_),
    .B1(_06405_),
    .B2(\reg_next_pc[23] ),
    .X(_06406_));
 sky130_fd_sc_hd__clkbuf_2 _27064_ (.A(_06406_),
    .X(_06407_));
 sky130_fd_sc_hd__a22o_1 _27065_ (.A1(_09750_),
    .A2(_06404_),
    .B1(_06391_),
    .B2(_06407_),
    .X(_00895_));
 sky130_fd_sc_hd__o22a_1 _27066_ (.A1(_10315_),
    .A2(_05201_),
    .B1(_06395_),
    .B2(\reg_next_pc[24] ),
    .X(_06408_));
 sky130_fd_sc_hd__and2_1 _27067_ (.A(_06394_),
    .B(_06408_),
    .X(_06409_));
 sky130_fd_sc_hd__clkbuf_2 _27068_ (.A(_06409_),
    .X(_06410_));
 sky130_fd_sc_hd__a22o_1 _27069_ (.A1(_09788_),
    .A2(_06404_),
    .B1(_06391_),
    .B2(_06410_),
    .X(_00896_));
 sky130_fd_sc_hd__clkbuf_2 _27070_ (.A(_06390_),
    .X(_06411_));
 sky130_fd_sc_hd__a22o_2 _27071_ (.A1(_10326_),
    .A2(_05210_),
    .B1(_06405_),
    .B2(\reg_next_pc[25] ),
    .X(_06412_));
 sky130_fd_sc_hd__clkbuf_2 _27072_ (.A(_06412_),
    .X(_06413_));
 sky130_fd_sc_hd__a22o_1 _27073_ (.A1(\reg_pc[25] ),
    .A2(_06404_),
    .B1(_06411_),
    .B2(_06413_),
    .X(_00897_));
 sky130_fd_sc_hd__o22a_1 _27074_ (.A1(_10315_),
    .A2(_05219_),
    .B1(_06395_),
    .B2(\reg_next_pc[26] ),
    .X(_06414_));
 sky130_fd_sc_hd__and2_1 _27075_ (.A(_06394_),
    .B(_06414_),
    .X(_06415_));
 sky130_fd_sc_hd__clkbuf_2 _27076_ (.A(_06415_),
    .X(_06416_));
 sky130_fd_sc_hd__a22o_1 _27077_ (.A1(_09894_),
    .A2(_06404_),
    .B1(_06411_),
    .B2(_06416_),
    .X(_00898_));
 sky130_fd_sc_hd__a22o_2 _27078_ (.A1(_10326_),
    .A2(_05227_),
    .B1(_06405_),
    .B2(\reg_next_pc[27] ),
    .X(_06417_));
 sky130_fd_sc_hd__clkbuf_2 _27079_ (.A(_06417_),
    .X(_06418_));
 sky130_fd_sc_hd__a22o_1 _27080_ (.A1(_09902_),
    .A2(_06404_),
    .B1(_06411_),
    .B2(_06418_),
    .X(_00899_));
 sky130_fd_sc_hd__o22a_1 _27081_ (.A1(_10315_),
    .A2(_05234_),
    .B1(_06395_),
    .B2(\reg_next_pc[28] ),
    .X(_06419_));
 sky130_fd_sc_hd__and2_1 _27082_ (.A(_06394_),
    .B(_06419_),
    .X(_06420_));
 sky130_fd_sc_hd__clkbuf_2 _27083_ (.A(_06420_),
    .X(_06421_));
 sky130_fd_sc_hd__a22o_1 _27084_ (.A1(\reg_pc[28] ),
    .A2(_06404_),
    .B1(_06411_),
    .B2(_06421_),
    .X(_00900_));
 sky130_fd_sc_hd__buf_2 _27085_ (.A(_06331_),
    .X(_06422_));
 sky130_fd_sc_hd__a22o_1 _27086_ (.A1(_10327_),
    .A2(_05242_),
    .B1(_06405_),
    .B2(\reg_next_pc[29] ),
    .X(_06423_));
 sky130_fd_sc_hd__clkbuf_2 _27087_ (.A(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__a22o_1 _27088_ (.A1(_09975_),
    .A2(_06422_),
    .B1(_06411_),
    .B2(_06424_),
    .X(_00901_));
 sky130_fd_sc_hd__o22a_1 _27089_ (.A1(_10315_),
    .A2(_05250_),
    .B1(_06395_),
    .B2(\reg_next_pc[30] ),
    .X(_06425_));
 sky130_fd_sc_hd__and2_1 _27090_ (.A(_06394_),
    .B(_06425_),
    .X(_06426_));
 sky130_fd_sc_hd__clkbuf_2 _27091_ (.A(_06426_),
    .X(_06427_));
 sky130_fd_sc_hd__a22o_1 _27092_ (.A1(\reg_pc[30] ),
    .A2(_06422_),
    .B1(_06411_),
    .B2(_06427_),
    .X(_00902_));
 sky130_fd_sc_hd__buf_2 _27093_ (.A(_06390_),
    .X(_06428_));
 sky130_fd_sc_hd__a22o_2 _27094_ (.A1(_10400_),
    .A2(_05258_),
    .B1(_06405_),
    .B2(\reg_next_pc[31] ),
    .X(_06429_));
 sky130_fd_sc_hd__a22o_1 _27095_ (.A1(\reg_pc[31] ),
    .A2(_06422_),
    .B1(_06428_),
    .B2(_06429_),
    .X(_00903_));
 sky130_fd_sc_hd__clkbuf_2 _27096_ (.A(_08307_),
    .X(_06430_));
 sky130_fd_sc_hd__clkbuf_2 _27097_ (.A(decoder_trigger),
    .X(_06431_));
 sky130_fd_sc_hd__nand2_2 _27098_ (.A(_08336_),
    .B(_06431_),
    .Y(_06432_));
 sky130_fd_sc_hd__buf_2 _27099_ (.A(_06432_),
    .X(_06433_));
 sky130_fd_sc_hd__or4_1 _27100_ (.A(_08207_),
    .B(_08547_),
    .C(_06430_),
    .D(_06433_),
    .X(_06434_));
 sky130_fd_sc_hd__xnor2_1 _27101_ (.A(_06337_),
    .B(_06434_),
    .Y(_06435_));
 sky130_fd_sc_hd__a22o_1 _27102_ (.A1(\reg_next_pc[1] ),
    .A2(_06422_),
    .B1(_06428_),
    .B2(_06435_),
    .X(_00904_));
 sky130_fd_sc_hd__buf_2 _27103_ (.A(_08176_),
    .X(_06436_));
 sky130_fd_sc_hd__or4_1 _27104_ (.A(\irq_pending[20] ),
    .B(\irq_pending[21] ),
    .C(\irq_pending[22] ),
    .D(\irq_pending[23] ),
    .X(_06437_));
 sky130_fd_sc_hd__or4_1 _27105_ (.A(\irq_pending[16] ),
    .B(\irq_pending[17] ),
    .C(\irq_pending[18] ),
    .D(\irq_pending[19] ),
    .X(_06438_));
 sky130_fd_sc_hd__nor2_1 _27106_ (.A(_06437_),
    .B(_06438_),
    .Y(_06439_));
 sky130_fd_sc_hd__or4_1 _27107_ (.A(\irq_pending[24] ),
    .B(\irq_pending[25] ),
    .C(\irq_pending[26] ),
    .D(\irq_pending[27] ),
    .X(_06440_));
 sky130_fd_sc_hd__or4_1 _27108_ (.A(\irq_pending[28] ),
    .B(\irq_pending[29] ),
    .C(\irq_pending[30] ),
    .D(\irq_pending[31] ),
    .X(_06441_));
 sky130_fd_sc_hd__nor2_1 _27109_ (.A(_06440_),
    .B(_06441_),
    .Y(_06442_));
 sky130_fd_sc_hd__or4_1 _27110_ (.A(\irq_pending[4] ),
    .B(\irq_pending[5] ),
    .C(\irq_pending[6] ),
    .D(\irq_pending[7] ),
    .X(_06443_));
 sky130_fd_sc_hd__or4_1 _27111_ (.A(\irq_pending[0] ),
    .B(\irq_pending[1] ),
    .C(\irq_pending[2] ),
    .D(\irq_pending[3] ),
    .X(_06444_));
 sky130_fd_sc_hd__nor2_1 _27112_ (.A(_06443_),
    .B(_06444_),
    .Y(_06445_));
 sky130_fd_sc_hd__or4_1 _27113_ (.A(\irq_pending[8] ),
    .B(\irq_pending[9] ),
    .C(\irq_pending[10] ),
    .D(\irq_pending[11] ),
    .X(_06446_));
 sky130_fd_sc_hd__or4_1 _27114_ (.A(\irq_pending[12] ),
    .B(\irq_pending[13] ),
    .C(\irq_pending[14] ),
    .D(\irq_pending[15] ),
    .X(_06447_));
 sky130_fd_sc_hd__nor2_1 _27115_ (.A(_06446_),
    .B(_06447_),
    .Y(_06448_));
 sky130_fd_sc_hd__nand4_4 _27116_ (.A(_06439_),
    .B(_06442_),
    .C(_06445_),
    .D(_06448_),
    .Y(_06449_));
 sky130_fd_sc_hd__nand2_2 _27117_ (.A(_08306_),
    .B(_06449_),
    .Y(_06450_));
 sky130_fd_sc_hd__nor2_2 _27118_ (.A(_08307_),
    .B(_06450_),
    .Y(_06451_));
 sky130_fd_sc_hd__or3b_1 _27119_ (.A(_06339_),
    .B(_06451_),
    .C_N(_08280_),
    .X(_06452_));
 sky130_fd_sc_hd__clkbuf_2 _27120_ (.A(_08336_),
    .X(_06453_));
 sky130_fd_sc_hd__buf_2 _27121_ (.A(_06453_),
    .X(_06454_));
 sky130_fd_sc_hd__clkbuf_4 _27122_ (.A(_06454_),
    .X(_06455_));
 sky130_fd_sc_hd__clkbuf_4 _27123_ (.A(_08303_),
    .X(_06456_));
 sky130_fd_sc_hd__and2_1 _27124_ (.A(\decoded_imm_uj[2] ),
    .B(_06338_),
    .X(_06457_));
 sky130_fd_sc_hd__or2_1 _27125_ (.A(\decoded_imm_uj[2] ),
    .B(_06338_),
    .X(_06458_));
 sky130_fd_sc_hd__and2b_1 _27126_ (.A_N(_06457_),
    .B(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__and3_1 _27127_ (.A(_08546_),
    .B(_06337_),
    .C(_06459_),
    .X(_06460_));
 sky130_fd_sc_hd__a21oi_1 _27128_ (.A1(_08546_),
    .A2(_06337_),
    .B1(_06459_),
    .Y(_06461_));
 sky130_fd_sc_hd__or3_1 _27129_ (.A(_06456_),
    .B(_06460_),
    .C(_06461_),
    .X(_06462_));
 sky130_fd_sc_hd__o21ai_1 _27130_ (.A1(_06455_),
    .A2(_06339_),
    .B1(_06462_),
    .Y(_06463_));
 sky130_fd_sc_hd__o2bb2a_1 _27131_ (.A1_N(_06339_),
    .A2_N(_06451_),
    .B1(_06463_),
    .B2(_08280_),
    .X(_06464_));
 sky130_fd_sc_hd__buf_2 _27132_ (.A(_06330_),
    .X(_06465_));
 sky130_fd_sc_hd__a32o_1 _27133_ (.A1(_06436_),
    .A2(_06452_),
    .A3(_06464_),
    .B1(_06465_),
    .B2(\reg_next_pc[2] ),
    .X(_00905_));
 sky130_fd_sc_hd__nor2_1 _27134_ (.A(_08277_),
    .B(_08278_),
    .Y(_06466_));
 sky130_fd_sc_hd__clkbuf_2 _27135_ (.A(_06466_),
    .X(_06467_));
 sky130_fd_sc_hd__clkbuf_2 _27136_ (.A(_08306_),
    .X(_06468_));
 sky130_fd_sc_hd__clkbuf_2 _27137_ (.A(_06449_),
    .X(_06469_));
 sky130_fd_sc_hd__and2_1 _27138_ (.A(_06338_),
    .B(_06342_),
    .X(_06470_));
 sky130_fd_sc_hd__nand2_1 _27139_ (.A(_06469_),
    .B(_06470_),
    .Y(_06471_));
 sky130_fd_sc_hd__a21o_1 _27140_ (.A1(_06339_),
    .A2(_06469_),
    .B1(_06342_),
    .X(_06472_));
 sky130_fd_sc_hd__clkbuf_4 _27141_ (.A(_08233_),
    .X(_06473_));
 sky130_fd_sc_hd__xor2_1 _27142_ (.A(\decoded_imm_uj[3] ),
    .B(_06341_),
    .X(_06474_));
 sky130_fd_sc_hd__a31o_1 _27143_ (.A1(\decoded_imm_uj[1] ),
    .A2(_06337_),
    .A3(_06458_),
    .B1(_06457_),
    .X(_06475_));
 sky130_fd_sc_hd__o21a_1 _27144_ (.A1(_06474_),
    .A2(_06475_),
    .B1(_08336_),
    .X(_06476_));
 sky130_fd_sc_hd__nand2_1 _27145_ (.A(_06474_),
    .B(_06475_),
    .Y(_06477_));
 sky130_fd_sc_hd__a2bb2o_1 _27146_ (.A1_N(_06453_),
    .A2_N(_06470_),
    .B1(_06476_),
    .B2(_06477_),
    .X(_06478_));
 sky130_fd_sc_hd__a211o_1 _27147_ (.A1(_06431_),
    .A2(_06339_),
    .B1(_06342_),
    .C1(_08304_),
    .X(_06479_));
 sky130_fd_sc_hd__o211a_1 _27148_ (.A1(_06473_),
    .A2(_06478_),
    .B1(_06479_),
    .C1(_08334_),
    .X(_06480_));
 sky130_fd_sc_hd__clkbuf_2 _27149_ (.A(_06430_),
    .X(_06481_));
 sky130_fd_sc_hd__a311o_1 _27150_ (.A1(_06468_),
    .A2(_06471_),
    .A3(_06472_),
    .B1(_06480_),
    .C1(_06481_),
    .X(_06482_));
 sky130_fd_sc_hd__o211a_1 _27151_ (.A1(_06467_),
    .A2(_06342_),
    .B1(_06482_),
    .C1(_06333_),
    .X(_06483_));
 sky130_fd_sc_hd__a21o_1 _27152_ (.A1(\reg_next_pc[3] ),
    .A2(_06332_),
    .B1(_06483_),
    .X(_00906_));
 sky130_fd_sc_hd__xnor2_1 _27153_ (.A(_06345_),
    .B(_06471_),
    .Y(_06484_));
 sky130_fd_sc_hd__nand2_2 _27154_ (.A(_06468_),
    .B(_06466_),
    .Y(_06485_));
 sky130_fd_sc_hd__clkbuf_2 _27155_ (.A(_06431_),
    .X(_06486_));
 sky130_fd_sc_hd__buf_2 _27156_ (.A(_06486_),
    .X(_06487_));
 sky130_fd_sc_hd__clkbuf_2 _27157_ (.A(_06431_),
    .X(_06488_));
 sky130_fd_sc_hd__and3_1 _27158_ (.A(_06338_),
    .B(_06342_),
    .C(_06344_),
    .X(_06489_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27159_ (.A(_06489_),
    .X(_06490_));
 sky130_fd_sc_hd__nand2_1 _27160_ (.A(_06488_),
    .B(_06490_),
    .Y(_06491_));
 sky130_fd_sc_hd__or2_1 _27161_ (.A(_06345_),
    .B(_06470_),
    .X(_06492_));
 sky130_fd_sc_hd__nand2_1 _27162_ (.A(\decoded_imm_uj[4] ),
    .B(_06345_),
    .Y(_06493_));
 sky130_fd_sc_hd__or2_1 _27163_ (.A(\decoded_imm_uj[4] ),
    .B(_06344_),
    .X(_06494_));
 sky130_fd_sc_hd__and2_1 _27164_ (.A(_06493_),
    .B(_06494_),
    .X(_06495_));
 sky130_fd_sc_hd__and2_1 _27165_ (.A(\decoded_imm_uj[3] ),
    .B(_06341_),
    .X(_06496_));
 sky130_fd_sc_hd__a21o_1 _27166_ (.A1(_06474_),
    .A2(_06475_),
    .B1(_06496_),
    .X(_06497_));
 sky130_fd_sc_hd__xor2_1 _27167_ (.A(_06495_),
    .B(_06497_),
    .X(_06498_));
 sky130_fd_sc_hd__a32o_1 _27168_ (.A1(_06433_),
    .A2(_06491_),
    .A3(_06492_),
    .B1(_06498_),
    .B2(_06454_),
    .X(_06499_));
 sky130_fd_sc_hd__o21ai_1 _27169_ (.A1(_06487_),
    .A2(_06345_),
    .B1(_06499_),
    .Y(_06500_));
 sky130_fd_sc_hd__nand2_1 _27170_ (.A(_08332_),
    .B(_06500_),
    .Y(_06501_));
 sky130_fd_sc_hd__o221a_1 _27171_ (.A1(_06467_),
    .A2(_06345_),
    .B1(_06484_),
    .B2(_06485_),
    .C1(_06501_),
    .X(_06502_));
 sky130_fd_sc_hd__a22o_1 _27172_ (.A1(\reg_next_pc[4] ),
    .A2(_06422_),
    .B1(_06428_),
    .B2(_06502_),
    .X(_00907_));
 sky130_fd_sc_hd__buf_2 _27173_ (.A(_06449_),
    .X(_06503_));
 sky130_fd_sc_hd__nand3_1 _27174_ (.A(_06349_),
    .B(_06503_),
    .C(_06490_),
    .Y(_06504_));
 sky130_fd_sc_hd__a21o_1 _27175_ (.A1(_06469_),
    .A2(_06490_),
    .B1(_06349_),
    .X(_06505_));
 sky130_fd_sc_hd__nand2_1 _27176_ (.A(_06348_),
    .B(_06490_),
    .Y(_06506_));
 sky130_fd_sc_hd__or2_1 _27177_ (.A(_06348_),
    .B(_06490_),
    .X(_06507_));
 sky130_fd_sc_hd__and2_1 _27178_ (.A(\decoded_imm_uj[5] ),
    .B(_06348_),
    .X(_06508_));
 sky130_fd_sc_hd__nor2_1 _27179_ (.A(\decoded_imm_uj[5] ),
    .B(_06348_),
    .Y(_06509_));
 sky130_fd_sc_hd__nor2_1 _27180_ (.A(_06508_),
    .B(_06509_),
    .Y(_06510_));
 sky130_fd_sc_hd__a21bo_1 _27181_ (.A1(_06494_),
    .A2(_06497_),
    .B1_N(_06493_),
    .X(_06511_));
 sky130_fd_sc_hd__and2_1 _27182_ (.A(_06510_),
    .B(_06511_),
    .X(_06512_));
 sky130_fd_sc_hd__o21ai_1 _27183_ (.A1(_06510_),
    .A2(_06511_),
    .B1(_08336_),
    .Y(_06513_));
 sky130_fd_sc_hd__nor2_1 _27184_ (.A(_06512_),
    .B(_06513_),
    .Y(_06514_));
 sky130_fd_sc_hd__a311o_1 _27185_ (.A1(_08303_),
    .A2(_06506_),
    .A3(_06507_),
    .B1(_06473_),
    .C1(_06514_),
    .X(_06515_));
 sky130_fd_sc_hd__o211a_1 _27186_ (.A1(_06486_),
    .A2(_06349_),
    .B1(_06515_),
    .C1(_08334_),
    .X(_06516_));
 sky130_fd_sc_hd__a311o_1 _27187_ (.A1(_06468_),
    .A2(_06504_),
    .A3(_06505_),
    .B1(_06516_),
    .C1(_06481_),
    .X(_06517_));
 sky130_fd_sc_hd__o211a_1 _27188_ (.A1(_06467_),
    .A2(_06349_),
    .B1(_06517_),
    .C1(_06333_),
    .X(_06518_));
 sky130_fd_sc_hd__a21o_1 _27189_ (.A1(\reg_next_pc[5] ),
    .A2(_06332_),
    .B1(_06518_),
    .X(_00908_));
 sky130_fd_sc_hd__or2_1 _27190_ (.A(\decoded_imm_uj[6] ),
    .B(_06352_),
    .X(_06519_));
 sky130_fd_sc_hd__nand2_1 _27191_ (.A(\decoded_imm_uj[6] ),
    .B(_06351_),
    .Y(_06520_));
 sky130_fd_sc_hd__nor2_1 _27192_ (.A(_06508_),
    .B(_06512_),
    .Y(_06521_));
 sky130_fd_sc_hd__a21oi_1 _27193_ (.A1(_06519_),
    .A2(_06520_),
    .B1(_06521_),
    .Y(_06522_));
 sky130_fd_sc_hd__a31o_1 _27194_ (.A1(_06521_),
    .A2(_06519_),
    .A3(_06520_),
    .B1(_06432_),
    .X(_06523_));
 sky130_fd_sc_hd__and3_1 _27195_ (.A(_06348_),
    .B(_06351_),
    .C(_06489_),
    .X(_06524_));
 sky130_fd_sc_hd__a21oi_1 _27196_ (.A1(_06349_),
    .A2(_06490_),
    .B1(_06352_),
    .Y(_06525_));
 sky130_fd_sc_hd__or2_1 _27197_ (.A(_06524_),
    .B(_06525_),
    .X(_06526_));
 sky130_fd_sc_hd__nand2_1 _27198_ (.A(_08338_),
    .B(_06526_),
    .Y(_06527_));
 sky130_fd_sc_hd__or2_1 _27199_ (.A(_06488_),
    .B(_06352_),
    .X(_06528_));
 sky130_fd_sc_hd__o211a_1 _27200_ (.A1(_06522_),
    .A2(_06523_),
    .B1(_06527_),
    .C1(_06528_),
    .X(_06529_));
 sky130_fd_sc_hd__and4_2 _27201_ (.A(_06439_),
    .B(_06442_),
    .C(_06445_),
    .D(_06448_),
    .X(_06530_));
 sky130_fd_sc_hd__nand2_1 _27202_ (.A(_08306_),
    .B(_06530_),
    .Y(_06531_));
 sky130_vsdinv _27203_ (.A(_06531_),
    .Y(_06532_));
 sky130_fd_sc_hd__a2bb2o_1 _27204_ (.A1_N(_06450_),
    .A2_N(_06526_),
    .B1(_06532_),
    .B2(_06352_),
    .X(_06533_));
 sky130_fd_sc_hd__buf_2 _27205_ (.A(_06430_),
    .X(_06534_));
 sky130_fd_sc_hd__a211o_1 _27206_ (.A1(_08334_),
    .A2(_06529_),
    .B1(_06533_),
    .C1(_06534_),
    .X(_06535_));
 sky130_fd_sc_hd__or2_1 _27207_ (.A(_06467_),
    .B(_06352_),
    .X(_06536_));
 sky130_fd_sc_hd__a32o_1 _27208_ (.A1(_06436_),
    .A2(_06535_),
    .A3(_06536_),
    .B1(_06465_),
    .B2(\reg_next_pc[6] ),
    .X(_00909_));
 sky130_vsdinv _27209_ (.A(_06355_),
    .Y(_06537_));
 sky130_fd_sc_hd__nand2_1 _27210_ (.A(_06355_),
    .B(_06524_),
    .Y(_06538_));
 sky130_fd_sc_hd__or2_1 _27211_ (.A(_06355_),
    .B(_06524_),
    .X(_06539_));
 sky130_fd_sc_hd__nand2_1 _27212_ (.A(_06538_),
    .B(_06539_),
    .Y(_06540_));
 sky130_fd_sc_hd__o221a_1 _27213_ (.A1(_06537_),
    .A2(_06531_),
    .B1(_06540_),
    .B2(_06450_),
    .C1(_06466_),
    .X(_06541_));
 sky130_fd_sc_hd__buf_2 _27214_ (.A(_06432_),
    .X(_06542_));
 sky130_fd_sc_hd__and2_1 _27215_ (.A(\decoded_imm_uj[7] ),
    .B(_06354_),
    .X(_06543_));
 sky130_fd_sc_hd__or2_1 _27216_ (.A(\decoded_imm_uj[7] ),
    .B(_06354_),
    .X(_06544_));
 sky130_fd_sc_hd__and2b_1 _27217_ (.A_N(_06543_),
    .B(_06544_),
    .X(_06545_));
 sky130_vsdinv _27218_ (.A(_06520_),
    .Y(_06546_));
 sky130_fd_sc_hd__a211o_1 _27219_ (.A1(_06510_),
    .A2(_06511_),
    .B1(_06546_),
    .C1(_06508_),
    .X(_06547_));
 sky130_fd_sc_hd__nand2_1 _27220_ (.A(_06519_),
    .B(_06547_),
    .Y(_06548_));
 sky130_fd_sc_hd__xnor2_1 _27221_ (.A(_06545_),
    .B(_06548_),
    .Y(_06549_));
 sky130_fd_sc_hd__a221oi_1 _27222_ (.A1(_06473_),
    .A2(_06537_),
    .B1(_06540_),
    .B2(_08338_),
    .C1(_06468_),
    .Y(_06550_));
 sky130_fd_sc_hd__o21ai_1 _27223_ (.A1(_06542_),
    .A2(_06549_),
    .B1(_06550_),
    .Y(_06551_));
 sky130_fd_sc_hd__o2bb2a_1 _27224_ (.A1_N(_06541_),
    .A2_N(_06551_),
    .B1(_06355_),
    .B2(_06467_),
    .X(_06552_));
 sky130_fd_sc_hd__a22o_1 _27225_ (.A1(\reg_next_pc[7] ),
    .A2(_06422_),
    .B1(_06428_),
    .B2(_06552_),
    .X(_00910_));
 sky130_fd_sc_hd__clkbuf_2 _27226_ (.A(_06331_),
    .X(_06553_));
 sky130_fd_sc_hd__xnor2_1 _27227_ (.A(_06358_),
    .B(_06538_),
    .Y(_06554_));
 sky130_fd_sc_hd__buf_2 _27228_ (.A(_06453_),
    .X(_06555_));
 sky130_fd_sc_hd__and2_1 _27229_ (.A(\decoded_imm_uj[8] ),
    .B(_06358_),
    .X(_06556_));
 sky130_fd_sc_hd__or2_1 _27230_ (.A(\decoded_imm_uj[8] ),
    .B(_06357_),
    .X(_06557_));
 sky130_fd_sc_hd__and2b_1 _27231_ (.A_N(_06556_),
    .B(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__a31o_1 _27232_ (.A1(_06519_),
    .A2(_06544_),
    .A3(_06547_),
    .B1(_06543_),
    .X(_06559_));
 sky130_fd_sc_hd__xnor2_1 _27233_ (.A(_06558_),
    .B(_06559_),
    .Y(_06560_));
 sky130_fd_sc_hd__a21oi_1 _27234_ (.A1(_06555_),
    .A2(_06560_),
    .B1(_08280_),
    .Y(_06561_));
 sky130_fd_sc_hd__o21a_1 _27235_ (.A1(_06555_),
    .A2(_06554_),
    .B1(_06561_),
    .X(_06562_));
 sky130_fd_sc_hd__or2_1 _27236_ (.A(_08307_),
    .B(_06450_),
    .X(_06563_));
 sky130_fd_sc_hd__and3_1 _27237_ (.A(_08280_),
    .B(_06358_),
    .C(_06563_),
    .X(_06564_));
 sky130_fd_sc_hd__a211o_1 _27238_ (.A1(_06451_),
    .A2(_06554_),
    .B1(_06562_),
    .C1(_06564_),
    .X(_06565_));
 sky130_fd_sc_hd__a22o_1 _27239_ (.A1(\reg_next_pc[8] ),
    .A2(_06553_),
    .B1(_06428_),
    .B2(_06565_),
    .X(_00911_));
 sky130_fd_sc_hd__and2_1 _27240_ (.A(\decoded_imm_uj[9] ),
    .B(_06360_),
    .X(_06566_));
 sky130_fd_sc_hd__nor2_1 _27241_ (.A(\decoded_imm_uj[9] ),
    .B(_06359_),
    .Y(_06567_));
 sky130_fd_sc_hd__nor2_1 _27242_ (.A(_06566_),
    .B(_06567_),
    .Y(_06568_));
 sky130_fd_sc_hd__a21o_1 _27243_ (.A1(_06557_),
    .A2(_06559_),
    .B1(_06556_),
    .X(_06569_));
 sky130_fd_sc_hd__and2_1 _27244_ (.A(_06568_),
    .B(_06569_),
    .X(_06570_));
 sky130_fd_sc_hd__o21ai_1 _27245_ (.A1(_06568_),
    .A2(_06569_),
    .B1(_06555_),
    .Y(_06571_));
 sky130_fd_sc_hd__or2b_1 _27246_ (.A(_06538_),
    .B_N(_06358_),
    .X(_06572_));
 sky130_fd_sc_hd__xor2_1 _27247_ (.A(_06360_),
    .B(_06572_),
    .X(_06573_));
 sky130_fd_sc_hd__clkbuf_2 _27248_ (.A(_06431_),
    .X(_06574_));
 sky130_fd_sc_hd__clkbuf_2 _27249_ (.A(_06574_),
    .X(_06575_));
 sky130_fd_sc_hd__o221a_1 _27250_ (.A1(_06570_),
    .A2(_06571_),
    .B1(_06573_),
    .B2(_06455_),
    .C1(_06575_),
    .X(_06576_));
 sky130_fd_sc_hd__o21ai_1 _27251_ (.A1(_06575_),
    .A2(_06360_),
    .B1(_08332_),
    .Y(_06577_));
 sky130_fd_sc_hd__buf_2 _27252_ (.A(_06466_),
    .X(_06578_));
 sky130_fd_sc_hd__nand2_1 _27253_ (.A(_06578_),
    .B(_06531_),
    .Y(_06579_));
 sky130_fd_sc_hd__o2bb2a_1 _27254_ (.A1_N(_06360_),
    .A2_N(_06579_),
    .B1(_06573_),
    .B2(_06563_),
    .X(_06580_));
 sky130_fd_sc_hd__o21ai_1 _27255_ (.A1(_06576_),
    .A2(_06577_),
    .B1(_06580_),
    .Y(_06581_));
 sky130_fd_sc_hd__a22o_1 _27256_ (.A1(\reg_next_pc[9] ),
    .A2(_06553_),
    .B1(_06428_),
    .B2(_06581_),
    .X(_00912_));
 sky130_fd_sc_hd__clkbuf_2 _27257_ (.A(decoder_trigger),
    .X(_06582_));
 sky130_fd_sc_hd__buf_2 _27258_ (.A(_06582_),
    .X(_06583_));
 sky130_fd_sc_hd__buf_2 _27259_ (.A(_06453_),
    .X(_06584_));
 sky130_fd_sc_hd__a21oi_1 _27260_ (.A1(_06557_),
    .A2(_06559_),
    .B1(_06556_),
    .Y(_06585_));
 sky130_fd_sc_hd__nand2_1 _27261_ (.A(\decoded_imm_uj[9] ),
    .B(_06359_),
    .Y(_06586_));
 sky130_fd_sc_hd__o21ai_1 _27262_ (.A1(_06567_),
    .A2(_06585_),
    .B1(_06586_),
    .Y(_06587_));
 sky130_fd_sc_hd__nor2_1 _27263_ (.A(\decoded_imm_uj[10] ),
    .B(_06365_),
    .Y(_06588_));
 sky130_fd_sc_hd__nand2_1 _27264_ (.A(\decoded_imm_uj[10] ),
    .B(_06364_),
    .Y(_06589_));
 sky130_fd_sc_hd__or2b_1 _27265_ (.A(_06588_),
    .B_N(_06589_),
    .X(_06590_));
 sky130_fd_sc_hd__xnor2_1 _27266_ (.A(_06587_),
    .B(_06590_),
    .Y(_06591_));
 sky130_fd_sc_hd__and3b_1 _27267_ (.A_N(_06572_),
    .B(_06359_),
    .C(_06363_),
    .X(_06592_));
 sky130_fd_sc_hd__a41o_1 _27268_ (.A1(_06355_),
    .A2(_06358_),
    .A3(_06360_),
    .A4(_06524_),
    .B1(_06365_),
    .X(_06593_));
 sky130_fd_sc_hd__or2b_1 _27269_ (.A(_06592_),
    .B_N(_06593_),
    .X(_06594_));
 sky130_fd_sc_hd__nand2_1 _27270_ (.A(_06582_),
    .B(_06594_),
    .Y(_06595_));
 sky130_fd_sc_hd__a22o_1 _27271_ (.A1(_06584_),
    .A2(_06591_),
    .B1(_06595_),
    .B2(_06432_),
    .X(_06596_));
 sky130_fd_sc_hd__o211a_1 _27272_ (.A1(_06583_),
    .A2(_06365_),
    .B1(_06596_),
    .C1(_08334_),
    .X(_06597_));
 sky130_fd_sc_hd__nor2_1 _27273_ (.A(_06450_),
    .B(_06594_),
    .Y(_06598_));
 sky130_fd_sc_hd__a2111o_1 _27274_ (.A1(_06365_),
    .A2(_06532_),
    .B1(_06597_),
    .C1(_06598_),
    .D1(_06534_),
    .X(_06599_));
 sky130_fd_sc_hd__or2_1 _27275_ (.A(_06578_),
    .B(_06365_),
    .X(_06600_));
 sky130_fd_sc_hd__a32o_1 _27276_ (.A1(_06436_),
    .A2(_06599_),
    .A3(_06600_),
    .B1(_06465_),
    .B2(\reg_next_pc[10] ),
    .X(_00913_));
 sky130_fd_sc_hd__buf_2 _27277_ (.A(_06390_),
    .X(_06601_));
 sky130_fd_sc_hd__nor2_1 _27278_ (.A(_08333_),
    .B(_08307_),
    .Y(_06602_));
 sky130_fd_sc_hd__clkbuf_2 _27279_ (.A(_06602_),
    .X(_06603_));
 sky130_fd_sc_hd__clkbuf_2 _27280_ (.A(_06603_),
    .X(_06604_));
 sky130_fd_sc_hd__buf_2 _27281_ (.A(_06503_),
    .X(_06605_));
 sky130_fd_sc_hd__xnor2_1 _27282_ (.A(_06368_),
    .B(_06592_),
    .Y(_06606_));
 sky130_fd_sc_hd__nand2_1 _27283_ (.A(_06605_),
    .B(_06606_),
    .Y(_06607_));
 sky130_fd_sc_hd__clkbuf_2 _27284_ (.A(_06449_),
    .X(_06608_));
 sky130_fd_sc_hd__or2_1 _27285_ (.A(_06368_),
    .B(_06608_),
    .X(_06609_));
 sky130_fd_sc_hd__and2_1 _27286_ (.A(_08554_),
    .B(_06367_),
    .X(_06610_));
 sky130_fd_sc_hd__nor2_1 _27287_ (.A(\decoded_imm_uj[11] ),
    .B(_06367_),
    .Y(_06611_));
 sky130_fd_sc_hd__nor2_1 _27288_ (.A(_06610_),
    .B(_06611_),
    .Y(_06612_));
 sky130_fd_sc_hd__o211a_1 _27289_ (.A1(_06567_),
    .A2(_06585_),
    .B1(_06589_),
    .C1(_06586_),
    .X(_06613_));
 sky130_fd_sc_hd__or2_1 _27290_ (.A(_06588_),
    .B(_06613_),
    .X(_06614_));
 sky130_fd_sc_hd__xnor2_1 _27291_ (.A(_06612_),
    .B(_06614_),
    .Y(_06615_));
 sky130_fd_sc_hd__nand2_1 _27292_ (.A(_08337_),
    .B(_06606_),
    .Y(_06616_));
 sky130_fd_sc_hd__o221a_1 _27293_ (.A1(_06486_),
    .A2(_06368_),
    .B1(_06615_),
    .B2(_06432_),
    .C1(_06616_),
    .X(_06617_));
 sky130_fd_sc_hd__a22o_1 _27294_ (.A1(_06481_),
    .A2(_06368_),
    .B1(_06617_),
    .B2(_08309_),
    .X(_06618_));
 sky130_fd_sc_hd__a31o_1 _27295_ (.A1(_06604_),
    .A2(_06607_),
    .A3(_06609_),
    .B1(_06618_),
    .X(_06619_));
 sky130_fd_sc_hd__a22o_1 _27296_ (.A1(\reg_next_pc[11] ),
    .A2(_06553_),
    .B1(_06601_),
    .B2(_06619_),
    .X(_00914_));
 sky130_fd_sc_hd__buf_2 _27297_ (.A(_06430_),
    .X(_06620_));
 sky130_fd_sc_hd__nand3_1 _27298_ (.A(_06367_),
    .B(_06369_),
    .C(_06592_),
    .Y(_06621_));
 sky130_fd_sc_hd__a21o_1 _27299_ (.A1(_06368_),
    .A2(_06592_),
    .B1(_06371_),
    .X(_06622_));
 sky130_fd_sc_hd__nand2_1 _27300_ (.A(_06621_),
    .B(_06622_),
    .Y(_06623_));
 sky130_vsdinv _27301_ (.A(_06623_),
    .Y(_06624_));
 sky130_fd_sc_hd__mux2_1 _27302_ (.A0(_06371_),
    .A1(_06624_),
    .S(_06608_),
    .X(_06625_));
 sky130_fd_sc_hd__nand2_1 _27303_ (.A(_08554_),
    .B(_06367_),
    .Y(_06626_));
 sky130_fd_sc_hd__o31a_1 _27304_ (.A1(_06588_),
    .A2(_06611_),
    .A3(_06613_),
    .B1(_06626_),
    .X(_06627_));
 sky130_fd_sc_hd__or2_1 _27305_ (.A(\decoded_imm_uj[12] ),
    .B(_06371_),
    .X(_06628_));
 sky130_fd_sc_hd__nand2_1 _27306_ (.A(\decoded_imm_uj[12] ),
    .B(_06370_),
    .Y(_06629_));
 sky130_fd_sc_hd__nand2_1 _27307_ (.A(_06628_),
    .B(_06629_),
    .Y(_06630_));
 sky130_fd_sc_hd__xor2_1 _27308_ (.A(_06627_),
    .B(_06630_),
    .X(_06631_));
 sky130_fd_sc_hd__nand2_2 _27309_ (.A(_06456_),
    .B(_06431_),
    .Y(_06632_));
 sky130_fd_sc_hd__o221a_1 _27310_ (.A1(_06486_),
    .A2(_06371_),
    .B1(_06624_),
    .B2(_06632_),
    .C1(_08308_),
    .X(_06633_));
 sky130_fd_sc_hd__o21a_1 _27311_ (.A1(_06542_),
    .A2(_06631_),
    .B1(_06633_),
    .X(_06634_));
 sky130_fd_sc_hd__a221o_1 _27312_ (.A1(_06620_),
    .A2(_06371_),
    .B1(_06625_),
    .B2(_06604_),
    .C1(_06634_),
    .X(_06635_));
 sky130_fd_sc_hd__a22o_1 _27313_ (.A1(\reg_next_pc[12] ),
    .A2(_06553_),
    .B1(_06601_),
    .B2(_06635_),
    .X(_00915_));
 sky130_fd_sc_hd__and2b_1 _27314_ (.A_N(_06621_),
    .B(_06374_),
    .X(_06636_));
 sky130_fd_sc_hd__and2b_1 _27315_ (.A_N(_06375_),
    .B(_06621_),
    .X(_06637_));
 sky130_fd_sc_hd__nor2_1 _27316_ (.A(_06636_),
    .B(_06637_),
    .Y(_06638_));
 sky130_fd_sc_hd__mux2_1 _27317_ (.A0(_06375_),
    .A1(_06638_),
    .S(_06503_),
    .X(_06639_));
 sky130_fd_sc_hd__and2_1 _27318_ (.A(\decoded_imm_uj[13] ),
    .B(_06375_),
    .X(_06640_));
 sky130_fd_sc_hd__or2_1 _27319_ (.A(\decoded_imm_uj[13] ),
    .B(_06374_),
    .X(_06641_));
 sky130_fd_sc_hd__and2b_1 _27320_ (.A_N(_06640_),
    .B(_06641_),
    .X(_06642_));
 sky130_fd_sc_hd__nand2_1 _27321_ (.A(_06627_),
    .B(_06629_),
    .Y(_06643_));
 sky130_fd_sc_hd__nand2_1 _27322_ (.A(_06628_),
    .B(_06643_),
    .Y(_06644_));
 sky130_fd_sc_hd__xnor2_1 _27323_ (.A(_06642_),
    .B(_06644_),
    .Y(_06645_));
 sky130_fd_sc_hd__o221a_1 _27324_ (.A1(_06486_),
    .A2(_06375_),
    .B1(_06638_),
    .B2(_06632_),
    .C1(_08308_),
    .X(_06646_));
 sky130_fd_sc_hd__o21a_1 _27325_ (.A1(_06542_),
    .A2(_06645_),
    .B1(_06646_),
    .X(_06647_));
 sky130_fd_sc_hd__a221o_1 _27326_ (.A1(_06620_),
    .A2(_06375_),
    .B1(_06639_),
    .B2(_06604_),
    .C1(_06647_),
    .X(_06648_));
 sky130_fd_sc_hd__a22o_1 _27327_ (.A1(\reg_next_pc[13] ),
    .A2(_06553_),
    .B1(_06601_),
    .B2(_06648_),
    .X(_00916_));
 sky130_fd_sc_hd__and2_1 _27328_ (.A(_06376_),
    .B(_06636_),
    .X(_06649_));
 sky130_fd_sc_hd__o21ba_1 _27329_ (.A1(_06378_),
    .A2(_06636_),
    .B1_N(_06649_),
    .X(_06650_));
 sky130_fd_sc_hd__mux2_1 _27330_ (.A0(_06378_),
    .A1(_06650_),
    .S(_06469_),
    .X(_06651_));
 sky130_fd_sc_hd__a31o_1 _27331_ (.A1(_06628_),
    .A2(_06641_),
    .A3(_06643_),
    .B1(_06640_),
    .X(_06652_));
 sky130_fd_sc_hd__or2_1 _27332_ (.A(\decoded_imm_uj[14] ),
    .B(_06377_),
    .X(_06653_));
 sky130_fd_sc_hd__nand2_1 _27333_ (.A(\decoded_imm_uj[14] ),
    .B(_06378_),
    .Y(_06654_));
 sky130_fd_sc_hd__nand2_1 _27334_ (.A(_06653_),
    .B(_06654_),
    .Y(_06655_));
 sky130_fd_sc_hd__xnor2_1 _27335_ (.A(_06652_),
    .B(_06655_),
    .Y(_06656_));
 sky130_fd_sc_hd__o221a_1 _27336_ (.A1(_06488_),
    .A2(_06378_),
    .B1(_06650_),
    .B2(_06632_),
    .C1(_08333_),
    .X(_06657_));
 sky130_fd_sc_hd__o21a_1 _27337_ (.A1(_06433_),
    .A2(_06656_),
    .B1(_06657_),
    .X(_06658_));
 sky130_fd_sc_hd__a211o_1 _27338_ (.A1(_06468_),
    .A2(_06651_),
    .B1(_06658_),
    .C1(_06534_),
    .X(_06659_));
 sky130_fd_sc_hd__or2_1 _27339_ (.A(_06578_),
    .B(_06378_),
    .X(_06660_));
 sky130_fd_sc_hd__a32o_1 _27340_ (.A1(_06436_),
    .A2(_06659_),
    .A3(_06660_),
    .B1(_06465_),
    .B2(\reg_next_pc[14] ),
    .X(_00917_));
 sky130_fd_sc_hd__and2_1 _27341_ (.A(\decoded_imm_uj[15] ),
    .B(_06379_),
    .X(_06661_));
 sky130_fd_sc_hd__nor2_1 _27342_ (.A(\decoded_imm_uj[15] ),
    .B(_06379_),
    .Y(_06662_));
 sky130_fd_sc_hd__nor2_1 _27343_ (.A(_06661_),
    .B(_06662_),
    .Y(_06663_));
 sky130_fd_sc_hd__a21bo_1 _27344_ (.A1(_06652_),
    .A2(_06653_),
    .B1_N(_06654_),
    .X(_06664_));
 sky130_fd_sc_hd__and2_1 _27345_ (.A(_06663_),
    .B(_06664_),
    .X(_06665_));
 sky130_fd_sc_hd__or2_1 _27346_ (.A(_06663_),
    .B(_06664_),
    .X(_06666_));
 sky130_fd_sc_hd__and3b_1 _27347_ (.A_N(_06665_),
    .B(_06453_),
    .C(_06666_),
    .X(_06667_));
 sky130_fd_sc_hd__xnor2_1 _27348_ (.A(_06380_),
    .B(_06649_),
    .Y(_06668_));
 sky130_fd_sc_hd__o21ai_1 _27349_ (.A1(_06584_),
    .A2(_06668_),
    .B1(_06488_),
    .Y(_06669_));
 sky130_fd_sc_hd__o221a_1 _27350_ (.A1(_06574_),
    .A2(_06380_),
    .B1(_06667_),
    .B2(_06669_),
    .C1(_08334_),
    .X(_06670_));
 sky130_fd_sc_hd__a2bb2o_1 _27351_ (.A1_N(_06450_),
    .A2_N(_06668_),
    .B1(_06532_),
    .B2(_06380_),
    .X(_06671_));
 sky130_fd_sc_hd__or3_1 _27352_ (.A(_06481_),
    .B(_06670_),
    .C(_06671_),
    .X(_06672_));
 sky130_fd_sc_hd__or2_1 _27353_ (.A(_06578_),
    .B(_06380_),
    .X(_06673_));
 sky130_fd_sc_hd__a32o_1 _27354_ (.A1(_06436_),
    .A2(_06672_),
    .A3(_06673_),
    .B1(_06346_),
    .B2(\reg_next_pc[15] ),
    .X(_00918_));
 sky130_fd_sc_hd__nand2_1 _27355_ (.A(\decoded_imm_uj[16] ),
    .B(_06382_),
    .Y(_06674_));
 sky130_fd_sc_hd__or2_1 _27356_ (.A(\decoded_imm_uj[16] ),
    .B(_06383_),
    .X(_06675_));
 sky130_fd_sc_hd__nand2_1 _27357_ (.A(_06674_),
    .B(_06675_),
    .Y(_06676_));
 sky130_fd_sc_hd__or2_1 _27358_ (.A(_06661_),
    .B(_06665_),
    .X(_06677_));
 sky130_fd_sc_hd__a21oi_1 _27359_ (.A1(_06676_),
    .A2(_06677_),
    .B1(_06542_),
    .Y(_06678_));
 sky130_fd_sc_hd__o21a_1 _27360_ (.A1(_06676_),
    .A2(_06677_),
    .B1(_06678_),
    .X(_06679_));
 sky130_fd_sc_hd__and3_1 _27361_ (.A(_06379_),
    .B(_06381_),
    .C(_06649_),
    .X(_06680_));
 sky130_fd_sc_hd__a21oi_1 _27362_ (.A1(_06380_),
    .A2(_06649_),
    .B1(_06383_),
    .Y(_06681_));
 sky130_fd_sc_hd__or2_1 _27363_ (.A(_06680_),
    .B(_06681_),
    .X(_06682_));
 sky130_fd_sc_hd__a2bb2o_1 _27364_ (.A1_N(_06575_),
    .A2_N(_06383_),
    .B1(_06682_),
    .B2(_08338_),
    .X(_06683_));
 sky130_fd_sc_hd__o21ai_1 _27365_ (.A1(_06679_),
    .A2(_06683_),
    .B1(_08332_),
    .Y(_06684_));
 sky130_fd_sc_hd__nor2_1 _27366_ (.A(_06530_),
    .B(_06682_),
    .Y(_06685_));
 sky130_fd_sc_hd__and2_1 _27367_ (.A(_06383_),
    .B(_06530_),
    .X(_06686_));
 sky130_fd_sc_hd__o32a_1 _27368_ (.A1(_06485_),
    .A2(_06685_),
    .A3(_06686_),
    .B1(_06383_),
    .B2(_06467_),
    .X(_06687_));
 sky130_fd_sc_hd__a32o_1 _27369_ (.A1(_06436_),
    .A2(_06684_),
    .A3(_06687_),
    .B1(_06346_),
    .B2(\reg_next_pc[16] ),
    .X(_00919_));
 sky130_fd_sc_hd__and2_1 _27370_ (.A(_06385_),
    .B(_06680_),
    .X(_06688_));
 sky130_fd_sc_hd__nor2_1 _27371_ (.A(_06386_),
    .B(_06680_),
    .Y(_06689_));
 sky130_fd_sc_hd__or2_1 _27372_ (.A(_06688_),
    .B(_06689_),
    .X(_06690_));
 sky130_fd_sc_hd__clkbuf_2 _27373_ (.A(_06469_),
    .X(_06691_));
 sky130_fd_sc_hd__nor2_1 _27374_ (.A(_06386_),
    .B(_06691_),
    .Y(_06692_));
 sky130_fd_sc_hd__a21oi_1 _27375_ (.A1(_06605_),
    .A2(_06690_),
    .B1(_06692_),
    .Y(_06693_));
 sky130_fd_sc_hd__nor2_1 _27376_ (.A(\decoded_imm_uj[17] ),
    .B(_06386_),
    .Y(_06694_));
 sky130_fd_sc_hd__and2_1 _27377_ (.A(\decoded_imm_uj[17] ),
    .B(_06385_),
    .X(_06695_));
 sky130_fd_sc_hd__nor2_1 _27378_ (.A(_06694_),
    .B(_06695_),
    .Y(_06696_));
 sky130_vsdinv _27379_ (.A(_06674_),
    .Y(_06697_));
 sky130_fd_sc_hd__a211o_1 _27380_ (.A1(_06675_),
    .A2(_06677_),
    .B1(_06696_),
    .C1(_06697_),
    .X(_06698_));
 sky130_fd_sc_hd__o311a_1 _27381_ (.A1(_06661_),
    .A2(_06665_),
    .A3(_06697_),
    .B1(_06675_),
    .C1(_06696_),
    .X(_06699_));
 sky130_fd_sc_hd__nor2_1 _27382_ (.A(_06456_),
    .B(_06699_),
    .Y(_06700_));
 sky130_fd_sc_hd__buf_2 _27383_ (.A(_08336_),
    .X(_06701_));
 sky130_fd_sc_hd__nor2_1 _27384_ (.A(_06701_),
    .B(_06690_),
    .Y(_06702_));
 sky130_fd_sc_hd__a211o_1 _27385_ (.A1(_06698_),
    .A2(_06700_),
    .B1(_06702_),
    .C1(_06473_),
    .X(_06703_));
 sky130_fd_sc_hd__o211a_1 _27386_ (.A1(_06487_),
    .A2(_06386_),
    .B1(_06703_),
    .C1(_08309_),
    .X(_06704_));
 sky130_fd_sc_hd__a221o_1 _27387_ (.A1(_06620_),
    .A2(_06386_),
    .B1(_06693_),
    .B2(_06604_),
    .C1(_06704_),
    .X(_06705_));
 sky130_fd_sc_hd__a22o_1 _27388_ (.A1(\reg_next_pc[17] ),
    .A2(_06553_),
    .B1(_06601_),
    .B2(_06705_),
    .X(_00920_));
 sky130_fd_sc_hd__clkbuf_2 _27389_ (.A(_06331_),
    .X(_06706_));
 sky130_fd_sc_hd__nand2_1 _27390_ (.A(\decoded_imm_uj[18] ),
    .B(_06388_),
    .Y(_06707_));
 sky130_fd_sc_hd__or2_1 _27391_ (.A(\decoded_imm_uj[18] ),
    .B(_06389_),
    .X(_06708_));
 sky130_fd_sc_hd__nor2_1 _27392_ (.A(_06695_),
    .B(_06699_),
    .Y(_06709_));
 sky130_fd_sc_hd__a21oi_1 _27393_ (.A1(_06707_),
    .A2(_06708_),
    .B1(_06709_),
    .Y(_06710_));
 sky130_fd_sc_hd__a31o_1 _27394_ (.A1(_06707_),
    .A2(_06708_),
    .A3(_06709_),
    .B1(_06433_),
    .X(_06711_));
 sky130_fd_sc_hd__nand2_1 _27395_ (.A(_06387_),
    .B(_06688_),
    .Y(_06712_));
 sky130_fd_sc_hd__o21ai_1 _27396_ (.A1(_06389_),
    .A2(_06688_),
    .B1(_06712_),
    .Y(_06713_));
 sky130_fd_sc_hd__o2bb2a_1 _27397_ (.A1_N(_08338_),
    .A2_N(_06713_),
    .B1(_06389_),
    .B2(_06488_),
    .X(_06714_));
 sky130_fd_sc_hd__o21a_1 _27398_ (.A1(_06710_),
    .A2(_06711_),
    .B1(_06714_),
    .X(_06715_));
 sky130_fd_sc_hd__nor2_1 _27399_ (.A(_06530_),
    .B(_06713_),
    .Y(_06716_));
 sky130_fd_sc_hd__a211o_1 _27400_ (.A1(_06389_),
    .A2(_06530_),
    .B1(_06716_),
    .C1(_06485_),
    .X(_06717_));
 sky130_fd_sc_hd__or2_1 _27401_ (.A(_06578_),
    .B(_06389_),
    .X(_06718_));
 sky130_fd_sc_hd__o311a_1 _27402_ (.A1(_06468_),
    .A2(_06534_),
    .A3(_06715_),
    .B1(_06717_),
    .C1(_06718_),
    .X(_06719_));
 sky130_fd_sc_hd__a22o_1 _27403_ (.A1(\reg_next_pc[18] ),
    .A2(_06706_),
    .B1(_06601_),
    .B2(_06719_),
    .X(_00921_));
 sky130_fd_sc_hd__and3_1 _27404_ (.A(_06387_),
    .B(_06392_),
    .C(_06688_),
    .X(_06720_));
 sky130_fd_sc_hd__a21oi_1 _27405_ (.A1(_06387_),
    .A2(_06688_),
    .B1(_06393_),
    .Y(_06721_));
 sky130_fd_sc_hd__or2_1 _27406_ (.A(_06720_),
    .B(_06721_),
    .X(_06722_));
 sky130_fd_sc_hd__clkbuf_2 _27407_ (.A(_06469_),
    .X(_06723_));
 sky130_fd_sc_hd__nor2_1 _27408_ (.A(_06393_),
    .B(_06723_),
    .Y(_06724_));
 sky130_fd_sc_hd__a21oi_1 _27409_ (.A1(_06605_),
    .A2(_06722_),
    .B1(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__clkbuf_4 _27410_ (.A(_06453_),
    .X(_06726_));
 sky130_fd_sc_hd__or2_1 _27411_ (.A(\decoded_imm_uj[19] ),
    .B(_06392_),
    .X(_06727_));
 sky130_fd_sc_hd__nand2_1 _27412_ (.A(\decoded_imm_uj[19] ),
    .B(_06393_),
    .Y(_06728_));
 sky130_fd_sc_hd__and2_1 _27413_ (.A(_06727_),
    .B(_06728_),
    .X(_06729_));
 sky130_vsdinv _27414_ (.A(_06707_),
    .Y(_06730_));
 sky130_fd_sc_hd__o31a_1 _27415_ (.A1(_06695_),
    .A2(_06699_),
    .A3(_06730_),
    .B1(_06708_),
    .X(_06731_));
 sky130_fd_sc_hd__or2_1 _27416_ (.A(_06729_),
    .B(_06731_),
    .X(_06732_));
 sky130_fd_sc_hd__o311ai_2 _27417_ (.A1(_06695_),
    .A2(_06699_),
    .A3(_06730_),
    .B1(_06708_),
    .C1(_06729_),
    .Y(_06733_));
 sky130_fd_sc_hd__o21ai_1 _27418_ (.A1(_06701_),
    .A2(_06722_),
    .B1(_06488_),
    .Y(_06734_));
 sky130_fd_sc_hd__a31o_1 _27419_ (.A1(_06726_),
    .A2(_06732_),
    .A3(_06733_),
    .B1(_06734_),
    .X(_06735_));
 sky130_fd_sc_hd__o211a_1 _27420_ (.A1(_06487_),
    .A2(_06393_),
    .B1(_06735_),
    .C1(_08309_),
    .X(_06736_));
 sky130_fd_sc_hd__a221o_1 _27421_ (.A1(_06620_),
    .A2(_06393_),
    .B1(_06725_),
    .B2(_06604_),
    .C1(_06736_),
    .X(_06737_));
 sky130_fd_sc_hd__a22o_1 _27422_ (.A1(\reg_next_pc[19] ),
    .A2(_06706_),
    .B1(_06601_),
    .B2(_06737_),
    .X(_00922_));
 sky130_fd_sc_hd__clkbuf_2 _27423_ (.A(_06390_),
    .X(_06738_));
 sky130_fd_sc_hd__clkbuf_2 _27424_ (.A(_06430_),
    .X(_06739_));
 sky130_fd_sc_hd__and2_1 _27425_ (.A(_06396_),
    .B(_06720_),
    .X(_06740_));
 sky130_fd_sc_hd__o21bai_1 _27426_ (.A1(_06398_),
    .A2(_06720_),
    .B1_N(_06740_),
    .Y(_06741_));
 sky130_vsdinv _27427_ (.A(_06741_),
    .Y(_06742_));
 sky130_fd_sc_hd__mux2_1 _27428_ (.A0(_06398_),
    .A1(_06742_),
    .S(_06503_),
    .X(_06743_));
 sky130_fd_sc_hd__clkbuf_2 _27429_ (.A(_06602_),
    .X(_06744_));
 sky130_fd_sc_hd__or2_1 _27430_ (.A(\decoded_imm_uj[20] ),
    .B(_06397_),
    .X(_06745_));
 sky130_fd_sc_hd__nand2_1 _27431_ (.A(\decoded_imm_uj[20] ),
    .B(_06398_),
    .Y(_06746_));
 sky130_fd_sc_hd__nand2_1 _27432_ (.A(_06745_),
    .B(_06746_),
    .Y(_06747_));
 sky130_fd_sc_hd__and2_1 _27433_ (.A(_06728_),
    .B(_06733_),
    .X(_06748_));
 sky130_fd_sc_hd__o21ai_1 _27434_ (.A1(_06747_),
    .A2(_06748_),
    .B1(_06584_),
    .Y(_06749_));
 sky130_fd_sc_hd__a21oi_1 _27435_ (.A1(_06747_),
    .A2(_06748_),
    .B1(_06749_),
    .Y(_06750_));
 sky130_fd_sc_hd__o21ai_1 _27436_ (.A1(_06454_),
    .A2(_06741_),
    .B1(_06574_),
    .Y(_06751_));
 sky130_fd_sc_hd__o221a_1 _27437_ (.A1(_06583_),
    .A2(_06398_),
    .B1(_06750_),
    .B2(_06751_),
    .C1(_08331_),
    .X(_06752_));
 sky130_fd_sc_hd__a221o_1 _27438_ (.A1(_06739_),
    .A2(_06398_),
    .B1(_06743_),
    .B2(_06744_),
    .C1(_06752_),
    .X(_06753_));
 sky130_fd_sc_hd__a22o_1 _27439_ (.A1(\reg_next_pc[20] ),
    .A2(_06706_),
    .B1(_06738_),
    .B2(_06753_),
    .X(_00923_));
 sky130_fd_sc_hd__xnor2_1 _27440_ (.A(_06399_),
    .B(_06740_),
    .Y(_06754_));
 sky130_fd_sc_hd__nor2_1 _27441_ (.A(_06400_),
    .B(_06723_),
    .Y(_06755_));
 sky130_fd_sc_hd__a21oi_1 _27442_ (.A1(_06605_),
    .A2(_06754_),
    .B1(_06755_),
    .Y(_06756_));
 sky130_fd_sc_hd__xor2_1 _27443_ (.A(\decoded_imm_uj[20] ),
    .B(_06399_),
    .X(_06757_));
 sky130_vsdinv _27444_ (.A(_06745_),
    .Y(_06758_));
 sky130_fd_sc_hd__a21oi_1 _27445_ (.A1(_06746_),
    .A2(_06748_),
    .B1(_06758_),
    .Y(_06759_));
 sky130_fd_sc_hd__or2_1 _27446_ (.A(_06757_),
    .B(_06759_),
    .X(_06760_));
 sky130_vsdinv _27447_ (.A(_06757_),
    .Y(_06761_));
 sky130_fd_sc_hd__a311o_1 _27448_ (.A1(_06728_),
    .A2(_06733_),
    .A3(_06746_),
    .B1(_06761_),
    .C1(_06758_),
    .X(_06762_));
 sky130_fd_sc_hd__o21ai_1 _27449_ (.A1(_06701_),
    .A2(_06754_),
    .B1(_06582_),
    .Y(_06763_));
 sky130_fd_sc_hd__a31o_1 _27450_ (.A1(_06726_),
    .A2(_06760_),
    .A3(_06762_),
    .B1(_06763_),
    .X(_06764_));
 sky130_fd_sc_hd__o211a_1 _27451_ (.A1(_06487_),
    .A2(_06400_),
    .B1(_06764_),
    .C1(_08309_),
    .X(_06765_));
 sky130_fd_sc_hd__a221o_1 _27452_ (.A1(_06739_),
    .A2(_06400_),
    .B1(_06756_),
    .B2(_06744_),
    .C1(_06765_),
    .X(_06766_));
 sky130_fd_sc_hd__a22o_1 _27453_ (.A1(\reg_next_pc[21] ),
    .A2(_06706_),
    .B1(_06738_),
    .B2(_06766_),
    .X(_00924_));
 sky130_fd_sc_hd__and3_1 _27454_ (.A(_06399_),
    .B(_06401_),
    .C(_06740_),
    .X(_06767_));
 sky130_fd_sc_hd__a21oi_1 _27455_ (.A1(_06400_),
    .A2(_06740_),
    .B1(_06403_),
    .Y(_06768_));
 sky130_fd_sc_hd__nor2_1 _27456_ (.A(_06767_),
    .B(_06768_),
    .Y(_06769_));
 sky130_fd_sc_hd__mux2_1 _27457_ (.A0(_06403_),
    .A1(_06769_),
    .S(_06503_),
    .X(_06770_));
 sky130_fd_sc_hd__xnor2_2 _27458_ (.A(\decoded_imm_uj[20] ),
    .B(_06402_),
    .Y(_06771_));
 sky130_fd_sc_hd__a21bo_1 _27459_ (.A1(_05552_),
    .A2(_06400_),
    .B1_N(_06762_),
    .X(_06772_));
 sky130_fd_sc_hd__nor2_1 _27460_ (.A(_06771_),
    .B(_06772_),
    .Y(_06773_));
 sky130_fd_sc_hd__a21o_1 _27461_ (.A1(_06771_),
    .A2(_06772_),
    .B1(_06433_),
    .X(_06774_));
 sky130_fd_sc_hd__o221a_1 _27462_ (.A1(_06486_),
    .A2(_06403_),
    .B1(_06769_),
    .B2(_06632_),
    .C1(_08308_),
    .X(_06775_));
 sky130_fd_sc_hd__o21a_1 _27463_ (.A1(_06773_),
    .A2(_06774_),
    .B1(_06775_),
    .X(_06776_));
 sky130_fd_sc_hd__a221o_1 _27464_ (.A1(_06739_),
    .A2(_06403_),
    .B1(_06770_),
    .B2(_06744_),
    .C1(_06776_),
    .X(_06777_));
 sky130_fd_sc_hd__a22o_1 _27465_ (.A1(\reg_next_pc[22] ),
    .A2(_06706_),
    .B1(_06738_),
    .B2(_06777_),
    .X(_00925_));
 sky130_fd_sc_hd__and2_1 _27466_ (.A(_06406_),
    .B(_06767_),
    .X(_06778_));
 sky130_fd_sc_hd__nor2_1 _27467_ (.A(_06407_),
    .B(_06767_),
    .Y(_06779_));
 sky130_fd_sc_hd__or2_1 _27468_ (.A(_06778_),
    .B(_06779_),
    .X(_06780_));
 sky130_fd_sc_hd__nor2_1 _27469_ (.A(_06407_),
    .B(_06723_),
    .Y(_06781_));
 sky130_fd_sc_hd__a21oi_1 _27470_ (.A1(_06605_),
    .A2(_06780_),
    .B1(_06781_),
    .Y(_06782_));
 sky130_fd_sc_hd__xor2_1 _27471_ (.A(_05549_),
    .B(_06406_),
    .X(_06783_));
 sky130_fd_sc_hd__o21ai_1 _27472_ (.A1(_06399_),
    .A2(_06403_),
    .B1(_05549_),
    .Y(_06784_));
 sky130_fd_sc_hd__o21ai_1 _27473_ (.A1(_06762_),
    .A2(_06771_),
    .B1(_06784_),
    .Y(_06785_));
 sky130_fd_sc_hd__and2_1 _27474_ (.A(_06783_),
    .B(_06785_),
    .X(_06786_));
 sky130_fd_sc_hd__o21ai_1 _27475_ (.A1(_06783_),
    .A2(_06785_),
    .B1(_06584_),
    .Y(_06787_));
 sky130_fd_sc_hd__nor2_1 _27476_ (.A(_06786_),
    .B(_06787_),
    .Y(_06788_));
 sky130_fd_sc_hd__o21ai_1 _27477_ (.A1(_06454_),
    .A2(_06780_),
    .B1(_06574_),
    .Y(_06789_));
 sky130_fd_sc_hd__o221a_1 _27478_ (.A1(_06583_),
    .A2(_06407_),
    .B1(_06788_),
    .B2(_06789_),
    .C1(_08331_),
    .X(_06790_));
 sky130_fd_sc_hd__a221o_1 _27479_ (.A1(_06739_),
    .A2(_06407_),
    .B1(_06782_),
    .B2(_06744_),
    .C1(_06790_),
    .X(_06791_));
 sky130_fd_sc_hd__a22o_1 _27480_ (.A1(\reg_next_pc[23] ),
    .A2(_06706_),
    .B1(_06738_),
    .B2(_06791_),
    .X(_00926_));
 sky130_fd_sc_hd__clkbuf_2 _27481_ (.A(_06331_),
    .X(_06792_));
 sky130_fd_sc_hd__or2_1 _27482_ (.A(_06410_),
    .B(_06691_),
    .X(_06793_));
 sky130_fd_sc_hd__nand2_1 _27483_ (.A(_06408_),
    .B(_06778_),
    .Y(_06794_));
 sky130_fd_sc_hd__o21ai_1 _27484_ (.A1(_06410_),
    .A2(_06778_),
    .B1(_06794_),
    .Y(_06795_));
 sky130_fd_sc_hd__nand2_1 _27485_ (.A(_06608_),
    .B(_06795_),
    .Y(_06796_));
 sky130_fd_sc_hd__a22o_1 _27486_ (.A1(_06481_),
    .A2(_06410_),
    .B1(_06796_),
    .B2(_06603_),
    .X(_06797_));
 sky130_fd_sc_hd__xnor2_2 _27487_ (.A(_05549_),
    .B(_06409_),
    .Y(_06798_));
 sky130_fd_sc_hd__a21oi_1 _27488_ (.A1(_05552_),
    .A2(_06407_),
    .B1(_06786_),
    .Y(_06799_));
 sky130_fd_sc_hd__o21ai_1 _27489_ (.A1(_06798_),
    .A2(_06799_),
    .B1(_06726_),
    .Y(_06800_));
 sky130_fd_sc_hd__a21oi_1 _27490_ (.A1(_06798_),
    .A2(_06799_),
    .B1(_06800_),
    .Y(_06801_));
 sky130_fd_sc_hd__o21ai_1 _27491_ (.A1(_06555_),
    .A2(_06795_),
    .B1(_06583_),
    .Y(_06802_));
 sky130_fd_sc_hd__o221a_1 _27492_ (.A1(_06575_),
    .A2(_06410_),
    .B1(_06801_),
    .B2(_06802_),
    .C1(_08332_),
    .X(_06803_));
 sky130_fd_sc_hd__a21o_1 _27493_ (.A1(_06793_),
    .A2(_06797_),
    .B1(_06803_),
    .X(_06804_));
 sky130_fd_sc_hd__a22o_1 _27494_ (.A1(\reg_next_pc[24] ),
    .A2(_06792_),
    .B1(_06738_),
    .B2(_06804_),
    .X(_00927_));
 sky130_fd_sc_hd__and3_1 _27495_ (.A(_06408_),
    .B(_06412_),
    .C(_06778_),
    .X(_06805_));
 sky130_fd_sc_hd__a21oi_1 _27496_ (.A1(_06408_),
    .A2(_06778_),
    .B1(_06413_),
    .Y(_06806_));
 sky130_fd_sc_hd__or2_1 _27497_ (.A(_06805_),
    .B(_06806_),
    .X(_06807_));
 sky130_fd_sc_hd__nor2_1 _27498_ (.A(_06413_),
    .B(_06723_),
    .Y(_06808_));
 sky130_fd_sc_hd__a21oi_1 _27499_ (.A1(_06691_),
    .A2(_06807_),
    .B1(_06808_),
    .Y(_06809_));
 sky130_fd_sc_hd__or3b_1 _27500_ (.A(_06762_),
    .B(_06771_),
    .C_N(_06783_),
    .X(_06810_));
 sky130_fd_sc_hd__o21ai_1 _27501_ (.A1(_06406_),
    .A2(_06410_),
    .B1(_05549_),
    .Y(_06811_));
 sky130_fd_sc_hd__o211ai_2 _27502_ (.A1(_06798_),
    .A2(_06810_),
    .B1(_06811_),
    .C1(_06784_),
    .Y(_06812_));
 sky130_fd_sc_hd__xor2_1 _27503_ (.A(_05550_),
    .B(_06412_),
    .X(_06813_));
 sky130_fd_sc_hd__or2_1 _27504_ (.A(_06812_),
    .B(_06813_),
    .X(_06814_));
 sky130_fd_sc_hd__nand2_1 _27505_ (.A(_06812_),
    .B(_06813_),
    .Y(_06815_));
 sky130_fd_sc_hd__o21ai_1 _27506_ (.A1(_06701_),
    .A2(_06807_),
    .B1(_06582_),
    .Y(_06816_));
 sky130_fd_sc_hd__a31o_1 _27507_ (.A1(_06726_),
    .A2(_06814_),
    .A3(_06815_),
    .B1(_06816_),
    .X(_06817_));
 sky130_fd_sc_hd__o211a_1 _27508_ (.A1(_06487_),
    .A2(_06413_),
    .B1(_06817_),
    .C1(_08309_),
    .X(_06818_));
 sky130_fd_sc_hd__a221o_1 _27509_ (.A1(_06739_),
    .A2(_06413_),
    .B1(_06809_),
    .B2(_06744_),
    .C1(_06818_),
    .X(_06819_));
 sky130_fd_sc_hd__a22o_1 _27510_ (.A1(\reg_next_pc[25] ),
    .A2(_06792_),
    .B1(_06738_),
    .B2(_06819_),
    .X(_00928_));
 sky130_fd_sc_hd__clkbuf_2 _27511_ (.A(_06390_),
    .X(_06820_));
 sky130_fd_sc_hd__and2_1 _27512_ (.A(_06414_),
    .B(_06805_),
    .X(_06821_));
 sky130_fd_sc_hd__o21bai_1 _27513_ (.A1(_06416_),
    .A2(_06805_),
    .B1_N(_06821_),
    .Y(_06822_));
 sky130_vsdinv _27514_ (.A(_06822_),
    .Y(_06823_));
 sky130_fd_sc_hd__mux2_1 _27515_ (.A0(_06416_),
    .A1(_06823_),
    .S(_06503_),
    .X(_06824_));
 sky130_fd_sc_hd__xor2_1 _27516_ (.A(_05549_),
    .B(_06415_),
    .X(_06825_));
 sky130_fd_sc_hd__a21bo_1 _27517_ (.A1(_05551_),
    .A2(_06413_),
    .B1_N(_06815_),
    .X(_06826_));
 sky130_fd_sc_hd__o21ai_1 _27518_ (.A1(_06825_),
    .A2(_06826_),
    .B1(_06584_),
    .Y(_06827_));
 sky130_fd_sc_hd__a21oi_1 _27519_ (.A1(_06825_),
    .A2(_06826_),
    .B1(_06827_),
    .Y(_06828_));
 sky130_fd_sc_hd__o21ai_1 _27520_ (.A1(_06454_),
    .A2(_06822_),
    .B1(_06574_),
    .Y(_06829_));
 sky130_fd_sc_hd__o221a_1 _27521_ (.A1(_06583_),
    .A2(_06416_),
    .B1(_06828_),
    .B2(_06829_),
    .C1(_08331_),
    .X(_06830_));
 sky130_fd_sc_hd__a221o_1 _27522_ (.A1(_06739_),
    .A2(_06416_),
    .B1(_06824_),
    .B2(_06744_),
    .C1(_06830_),
    .X(_06831_));
 sky130_fd_sc_hd__a22o_1 _27523_ (.A1(\reg_next_pc[26] ),
    .A2(_06792_),
    .B1(_06820_),
    .B2(_06831_),
    .X(_00929_));
 sky130_fd_sc_hd__xnor2_1 _27524_ (.A(_06417_),
    .B(_06821_),
    .Y(_06832_));
 sky130_fd_sc_hd__nor2_1 _27525_ (.A(_06418_),
    .B(_06723_),
    .Y(_06833_));
 sky130_fd_sc_hd__a21oi_1 _27526_ (.A1(_06691_),
    .A2(_06832_),
    .B1(_06833_),
    .Y(_06834_));
 sky130_fd_sc_hd__xor2_1 _27527_ (.A(_05550_),
    .B(_06417_),
    .X(_06835_));
 sky130_fd_sc_hd__and3_1 _27528_ (.A(_06812_),
    .B(_06813_),
    .C(_06825_),
    .X(_06836_));
 sky130_fd_sc_hd__o21a_1 _27529_ (.A1(_06412_),
    .A2(_06416_),
    .B1(_05550_),
    .X(_06837_));
 sky130_fd_sc_hd__or2_1 _27530_ (.A(_06836_),
    .B(_06837_),
    .X(_06838_));
 sky130_fd_sc_hd__or2_1 _27531_ (.A(_06835_),
    .B(_06838_),
    .X(_06839_));
 sky130_fd_sc_hd__nand2_1 _27532_ (.A(_06835_),
    .B(_06838_),
    .Y(_06840_));
 sky130_fd_sc_hd__o21ai_1 _27533_ (.A1(_06701_),
    .A2(_06832_),
    .B1(_06582_),
    .Y(_06841_));
 sky130_fd_sc_hd__a31o_1 _27534_ (.A1(_06726_),
    .A2(_06839_),
    .A3(_06840_),
    .B1(_06841_),
    .X(_06842_));
 sky130_fd_sc_hd__o211a_1 _27535_ (.A1(_06487_),
    .A2(_06418_),
    .B1(_06842_),
    .C1(_08331_),
    .X(_06843_));
 sky130_fd_sc_hd__a221o_1 _27536_ (.A1(_06534_),
    .A2(_06418_),
    .B1(_06834_),
    .B2(_06603_),
    .C1(_06843_),
    .X(_06844_));
 sky130_fd_sc_hd__a22o_1 _27537_ (.A1(\reg_next_pc[27] ),
    .A2(_06792_),
    .B1(_06820_),
    .B2(_06844_),
    .X(_00930_));
 sky130_fd_sc_hd__and3_1 _27538_ (.A(_06417_),
    .B(_06419_),
    .C(_06821_),
    .X(_06845_));
 sky130_fd_sc_hd__a21oi_1 _27539_ (.A1(_06418_),
    .A2(_06821_),
    .B1(_06421_),
    .Y(_06846_));
 sky130_fd_sc_hd__or2_1 _27540_ (.A(_06845_),
    .B(_06846_),
    .X(_06847_));
 sky130_fd_sc_hd__xor2_1 _27541_ (.A(_05550_),
    .B(_06420_),
    .X(_06848_));
 sky130_fd_sc_hd__a21bo_1 _27542_ (.A1(_05552_),
    .A2(_06418_),
    .B1_N(_06840_),
    .X(_06849_));
 sky130_fd_sc_hd__nor2_1 _27543_ (.A(_06848_),
    .B(_06849_),
    .Y(_06850_));
 sky130_fd_sc_hd__a21o_1 _27544_ (.A1(_06848_),
    .A2(_06849_),
    .B1(_06456_),
    .X(_06851_));
 sky130_fd_sc_hd__o221a_1 _27545_ (.A1(_06455_),
    .A2(_06847_),
    .B1(_06850_),
    .B2(_06851_),
    .C1(_06575_),
    .X(_06852_));
 sky130_fd_sc_hd__o21ai_1 _27546_ (.A1(_06575_),
    .A2(_06421_),
    .B1(_08332_),
    .Y(_06853_));
 sky130_fd_sc_hd__nand2_1 _27547_ (.A(_06608_),
    .B(_06847_),
    .Y(_06854_));
 sky130_fd_sc_hd__a22o_1 _27548_ (.A1(_06481_),
    .A2(_06421_),
    .B1(_06854_),
    .B2(_06603_),
    .X(_06855_));
 sky130_fd_sc_hd__o21ai_1 _27549_ (.A1(_06421_),
    .A2(_06605_),
    .B1(_06855_),
    .Y(_06856_));
 sky130_fd_sc_hd__o21ai_1 _27550_ (.A1(_06852_),
    .A2(_06853_),
    .B1(_06856_),
    .Y(_06857_));
 sky130_fd_sc_hd__a22o_1 _27551_ (.A1(\reg_next_pc[28] ),
    .A2(_06792_),
    .B1(_06820_),
    .B2(_06857_),
    .X(_00931_));
 sky130_fd_sc_hd__and2_1 _27552_ (.A(_06423_),
    .B(_06845_),
    .X(_06858_));
 sky130_fd_sc_hd__nor2_1 _27553_ (.A(_06424_),
    .B(_06845_),
    .Y(_06859_));
 sky130_fd_sc_hd__or2_1 _27554_ (.A(_06858_),
    .B(_06859_),
    .X(_06860_));
 sky130_fd_sc_hd__nor2_1 _27555_ (.A(_06424_),
    .B(_06723_),
    .Y(_06861_));
 sky130_fd_sc_hd__a21oi_1 _27556_ (.A1(_06691_),
    .A2(_06860_),
    .B1(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__xor2_1 _27557_ (.A(_05551_),
    .B(_06423_),
    .X(_06863_));
 sky130_fd_sc_hd__o21a_1 _27558_ (.A1(_06417_),
    .A2(_06421_),
    .B1(_05550_),
    .X(_06864_));
 sky130_fd_sc_hd__a311o_1 _27559_ (.A1(_06835_),
    .A2(_06836_),
    .A3(_06848_),
    .B1(_06864_),
    .C1(_06837_),
    .X(_06865_));
 sky130_fd_sc_hd__or2_1 _27560_ (.A(_06863_),
    .B(_06865_),
    .X(_06866_));
 sky130_fd_sc_hd__nand2_1 _27561_ (.A(_06863_),
    .B(_06865_),
    .Y(_06867_));
 sky130_fd_sc_hd__o21ai_1 _27562_ (.A1(_06701_),
    .A2(_06860_),
    .B1(_06582_),
    .Y(_06868_));
 sky130_fd_sc_hd__a31o_1 _27563_ (.A1(_06584_),
    .A2(_06866_),
    .A3(_06867_),
    .B1(_06868_),
    .X(_06869_));
 sky130_fd_sc_hd__o211a_1 _27564_ (.A1(_06583_),
    .A2(_06424_),
    .B1(_06869_),
    .C1(_08331_),
    .X(_06870_));
 sky130_fd_sc_hd__a221o_1 _27565_ (.A1(_06534_),
    .A2(_06424_),
    .B1(_06862_),
    .B2(_06603_),
    .C1(_06870_),
    .X(_06871_));
 sky130_fd_sc_hd__a22o_1 _27566_ (.A1(\reg_next_pc[29] ),
    .A2(_06792_),
    .B1(_06820_),
    .B2(_06871_),
    .X(_00932_));
 sky130_fd_sc_hd__nand2_1 _27567_ (.A(_05551_),
    .B(_06426_),
    .Y(_06872_));
 sky130_vsdinv _27568_ (.A(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__nor2_1 _27569_ (.A(_05551_),
    .B(_06427_),
    .Y(_06874_));
 sky130_fd_sc_hd__nor2_1 _27570_ (.A(_06873_),
    .B(_06874_),
    .Y(_06875_));
 sky130_fd_sc_hd__a21boi_1 _27571_ (.A1(_05551_),
    .A2(_06424_),
    .B1_N(_06867_),
    .Y(_06876_));
 sky130_fd_sc_hd__xnor2_1 _27572_ (.A(_06875_),
    .B(_06876_),
    .Y(_06877_));
 sky130_fd_sc_hd__o21a_1 _27573_ (.A1(_06574_),
    .A2(_06427_),
    .B1(_08308_),
    .X(_06878_));
 sky130_fd_sc_hd__nand2_1 _27574_ (.A(_06425_),
    .B(_06858_),
    .Y(_06879_));
 sky130_fd_sc_hd__o21ai_1 _27575_ (.A1(_06427_),
    .A2(_06858_),
    .B1(_06879_),
    .Y(_06880_));
 sky130_fd_sc_hd__nand2_1 _27576_ (.A(_08338_),
    .B(_06880_),
    .Y(_06881_));
 sky130_fd_sc_hd__o211a_1 _27577_ (.A1(_06542_),
    .A2(_06877_),
    .B1(_06878_),
    .C1(_06881_),
    .X(_06882_));
 sky130_fd_sc_hd__nand2_1 _27578_ (.A(_06608_),
    .B(_06880_),
    .Y(_06883_));
 sky130_fd_sc_hd__o211a_1 _27579_ (.A1(_06427_),
    .A2(_06691_),
    .B1(_06883_),
    .C1(_06603_),
    .X(_06884_));
 sky130_fd_sc_hd__a211o_1 _27580_ (.A1(_06620_),
    .A2(_06427_),
    .B1(_06882_),
    .C1(_06884_),
    .X(_06885_));
 sky130_fd_sc_hd__a22o_1 _27581_ (.A1(\reg_next_pc[30] ),
    .A2(_06465_),
    .B1(_06820_),
    .B2(_06885_),
    .X(_00933_));
 sky130_fd_sc_hd__xnor2_1 _27582_ (.A(_06429_),
    .B(_06879_),
    .Y(_06886_));
 sky130_fd_sc_hd__mux2_1 _27583_ (.A0(_06429_),
    .A1(_06886_),
    .S(_06608_),
    .X(_06887_));
 sky130_fd_sc_hd__o211a_1 _27584_ (.A1(_06473_),
    .A2(_06430_),
    .B1(_06485_),
    .C1(_06429_),
    .X(_06888_));
 sky130_fd_sc_hd__a21oi_1 _27585_ (.A1(_06872_),
    .A2(_06876_),
    .B1(_06874_),
    .Y(_06889_));
 sky130_fd_sc_hd__xnor2_1 _27586_ (.A(_05552_),
    .B(_06429_),
    .Y(_06890_));
 sky130_fd_sc_hd__xnor2_1 _27587_ (.A(_06889_),
    .B(_06890_),
    .Y(_06891_));
 sky130_fd_sc_hd__o21ba_1 _27588_ (.A1(_06454_),
    .A2(_06886_),
    .B1_N(_08279_),
    .X(_06892_));
 sky130_fd_sc_hd__o21a_1 _27589_ (.A1(_06456_),
    .A2(_06891_),
    .B1(_06892_),
    .X(_06893_));
 sky130_fd_sc_hd__a211o_1 _27590_ (.A1(_06604_),
    .A2(_06887_),
    .B1(_06888_),
    .C1(_06893_),
    .X(_06894_));
 sky130_fd_sc_hd__a22o_1 _27591_ (.A1(\reg_next_pc[31] ),
    .A2(_06465_),
    .B1(_06820_),
    .B2(_06894_),
    .X(_00934_));
 sky130_fd_sc_hd__nor2_1 _27592_ (.A(_08655_),
    .B(_08521_),
    .Y(_00935_));
 sky130_fd_sc_hd__o21ai_1 _27593_ (.A1(_08655_),
    .A2(\count_cycle[1] ),
    .B1(_06180_),
    .Y(_06895_));
 sky130_fd_sc_hd__a21oi_1 _27594_ (.A1(_08655_),
    .A2(\count_cycle[1] ),
    .B1(_06895_),
    .Y(_00936_));
 sky130_fd_sc_hd__and3_1 _27595_ (.A(_08655_),
    .B(\count_cycle[1] ),
    .C(\count_cycle[2] ),
    .X(_06896_));
 sky130_fd_sc_hd__a21o_1 _27596_ (.A1(_08655_),
    .A2(\count_cycle[1] ),
    .B1(\count_cycle[2] ),
    .X(_06897_));
 sky130_fd_sc_hd__and3b_1 _27597_ (.A_N(_06896_),
    .B(_06302_),
    .C(_06897_),
    .X(_06898_));
 sky130_fd_sc_hd__clkbuf_1 _27598_ (.A(_06898_),
    .X(_00937_));
 sky130_fd_sc_hd__and4_2 _27599_ (.A(\count_cycle[0] ),
    .B(\count_cycle[1] ),
    .C(\count_cycle[2] ),
    .D(\count_cycle[3] ),
    .X(_06899_));
 sky130_fd_sc_hd__o21ai_1 _27600_ (.A1(\count_cycle[3] ),
    .A2(_06896_),
    .B1(_06324_),
    .Y(_06900_));
 sky130_fd_sc_hd__nor2_1 _27601_ (.A(_06899_),
    .B(_06900_),
    .Y(_00938_));
 sky130_fd_sc_hd__a21oi_1 _27602_ (.A1(\count_cycle[4] ),
    .A2(_06899_),
    .B1(_06286_),
    .Y(_06901_));
 sky130_fd_sc_hd__o21a_1 _27603_ (.A1(\count_cycle[4] ),
    .A2(_06899_),
    .B1(_06901_),
    .X(_00939_));
 sky130_fd_sc_hd__and3_1 _27604_ (.A(\count_cycle[4] ),
    .B(\count_cycle[5] ),
    .C(_06899_),
    .X(_06902_));
 sky130_fd_sc_hd__a21o_1 _27605_ (.A1(\count_cycle[4] ),
    .A2(_06899_),
    .B1(\count_cycle[5] ),
    .X(_06903_));
 sky130_fd_sc_hd__and3b_1 _27606_ (.A_N(_06902_),
    .B(_06302_),
    .C(_06903_),
    .X(_06904_));
 sky130_fd_sc_hd__clkbuf_1 _27607_ (.A(_06904_),
    .X(_00940_));
 sky130_fd_sc_hd__and4_2 _27608_ (.A(\count_cycle[4] ),
    .B(\count_cycle[5] ),
    .C(\count_cycle[6] ),
    .D(_06899_),
    .X(_06905_));
 sky130_fd_sc_hd__o21ai_1 _27609_ (.A1(\count_cycle[6] ),
    .A2(_06902_),
    .B1(_06324_),
    .Y(_06906_));
 sky130_fd_sc_hd__nor2_1 _27610_ (.A(_06905_),
    .B(_06906_),
    .Y(_00941_));
 sky130_fd_sc_hd__clkbuf_2 _27611_ (.A(_06200_),
    .X(_06907_));
 sky130_fd_sc_hd__a21oi_1 _27612_ (.A1(\count_cycle[7] ),
    .A2(_06905_),
    .B1(_06907_),
    .Y(_06908_));
 sky130_fd_sc_hd__o21a_1 _27613_ (.A1(\count_cycle[7] ),
    .A2(_06905_),
    .B1(_06908_),
    .X(_00942_));
 sky130_fd_sc_hd__and3_1 _27614_ (.A(\count_cycle[7] ),
    .B(\count_cycle[8] ),
    .C(_06905_),
    .X(_06909_));
 sky130_fd_sc_hd__a21o_1 _27615_ (.A1(\count_cycle[7] ),
    .A2(_06905_),
    .B1(\count_cycle[8] ),
    .X(_06910_));
 sky130_fd_sc_hd__and3b_1 _27616_ (.A_N(_06909_),
    .B(_06302_),
    .C(_06910_),
    .X(_06911_));
 sky130_fd_sc_hd__clkbuf_1 _27617_ (.A(_06911_),
    .X(_00943_));
 sky130_fd_sc_hd__and4_1 _27618_ (.A(\count_cycle[7] ),
    .B(\count_cycle[8] ),
    .C(\count_cycle[9] ),
    .D(_06905_),
    .X(_06912_));
 sky130_fd_sc_hd__o21ai_1 _27619_ (.A1(\count_cycle[9] ),
    .A2(_06909_),
    .B1(_06324_),
    .Y(_06913_));
 sky130_fd_sc_hd__nor2_1 _27620_ (.A(_06912_),
    .B(_06913_),
    .Y(_00944_));
 sky130_fd_sc_hd__a21oi_1 _27621_ (.A1(\count_cycle[10] ),
    .A2(_06912_),
    .B1(_06907_),
    .Y(_06914_));
 sky130_fd_sc_hd__o21a_1 _27622_ (.A1(\count_cycle[10] ),
    .A2(_06912_),
    .B1(_06914_),
    .X(_00945_));
 sky130_fd_sc_hd__and3_1 _27623_ (.A(\count_cycle[10] ),
    .B(\count_cycle[11] ),
    .C(_06912_),
    .X(_06915_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27624_ (.A(_08505_),
    .X(_06916_));
 sky130_fd_sc_hd__a21o_1 _27625_ (.A1(\count_cycle[10] ),
    .A2(_06912_),
    .B1(\count_cycle[11] ),
    .X(_06917_));
 sky130_fd_sc_hd__and3b_1 _27626_ (.A_N(_06915_),
    .B(_06916_),
    .C(_06917_),
    .X(_06918_));
 sky130_fd_sc_hd__clkbuf_1 _27627_ (.A(_06918_),
    .X(_00946_));
 sky130_fd_sc_hd__and4_2 _27628_ (.A(\count_cycle[10] ),
    .B(\count_cycle[11] ),
    .C(\count_cycle[12] ),
    .D(_06912_),
    .X(_06919_));
 sky130_fd_sc_hd__o21ai_1 _27629_ (.A1(\count_cycle[12] ),
    .A2(_06915_),
    .B1(_06324_),
    .Y(_06920_));
 sky130_fd_sc_hd__nor2_1 _27630_ (.A(_06919_),
    .B(_06920_),
    .Y(_00947_));
 sky130_fd_sc_hd__a21oi_1 _27631_ (.A1(\count_cycle[13] ),
    .A2(_06919_),
    .B1(_06907_),
    .Y(_06921_));
 sky130_fd_sc_hd__o21a_1 _27632_ (.A1(\count_cycle[13] ),
    .A2(_06919_),
    .B1(_06921_),
    .X(_00948_));
 sky130_fd_sc_hd__and3_1 _27633_ (.A(\count_cycle[13] ),
    .B(\count_cycle[14] ),
    .C(_06919_),
    .X(_06922_));
 sky130_fd_sc_hd__a21o_1 _27634_ (.A1(\count_cycle[13] ),
    .A2(_06919_),
    .B1(\count_cycle[14] ),
    .X(_06923_));
 sky130_fd_sc_hd__and3b_1 _27635_ (.A_N(_06922_),
    .B(_06916_),
    .C(_06923_),
    .X(_06924_));
 sky130_fd_sc_hd__clkbuf_1 _27636_ (.A(_06924_),
    .X(_00949_));
 sky130_fd_sc_hd__and4_1 _27637_ (.A(\count_cycle[13] ),
    .B(\count_cycle[14] ),
    .C(\count_cycle[15] ),
    .D(_06919_),
    .X(_06925_));
 sky130_fd_sc_hd__clkbuf_2 _27638_ (.A(_06235_),
    .X(_06926_));
 sky130_fd_sc_hd__o21ai_1 _27639_ (.A1(\count_cycle[15] ),
    .A2(_06922_),
    .B1(_06926_),
    .Y(_06927_));
 sky130_fd_sc_hd__nor2_1 _27640_ (.A(_06925_),
    .B(_06927_),
    .Y(_00950_));
 sky130_fd_sc_hd__a21oi_1 _27641_ (.A1(\count_cycle[16] ),
    .A2(_06925_),
    .B1(_06907_),
    .Y(_06928_));
 sky130_fd_sc_hd__o21a_1 _27642_ (.A1(\count_cycle[16] ),
    .A2(_06925_),
    .B1(_06928_),
    .X(_00951_));
 sky130_fd_sc_hd__and3_1 _27643_ (.A(\count_cycle[16] ),
    .B(\count_cycle[17] ),
    .C(_06925_),
    .X(_06929_));
 sky130_fd_sc_hd__a21o_1 _27644_ (.A1(\count_cycle[16] ),
    .A2(_06925_),
    .B1(\count_cycle[17] ),
    .X(_06930_));
 sky130_fd_sc_hd__and3b_1 _27645_ (.A_N(_06929_),
    .B(_06916_),
    .C(_06930_),
    .X(_06931_));
 sky130_fd_sc_hd__clkbuf_1 _27646_ (.A(_06931_),
    .X(_00952_));
 sky130_fd_sc_hd__and4_1 _27647_ (.A(\count_cycle[16] ),
    .B(\count_cycle[17] ),
    .C(\count_cycle[18] ),
    .D(_06925_),
    .X(_06932_));
 sky130_fd_sc_hd__o21ai_1 _27648_ (.A1(\count_cycle[18] ),
    .A2(_06929_),
    .B1(_06926_),
    .Y(_06933_));
 sky130_fd_sc_hd__nor2_1 _27649_ (.A(_06932_),
    .B(_06933_),
    .Y(_00953_));
 sky130_fd_sc_hd__a21oi_1 _27650_ (.A1(\count_cycle[19] ),
    .A2(_06932_),
    .B1(_06907_),
    .Y(_06934_));
 sky130_fd_sc_hd__o21a_1 _27651_ (.A1(\count_cycle[19] ),
    .A2(_06932_),
    .B1(_06934_),
    .X(_00954_));
 sky130_fd_sc_hd__and3_1 _27652_ (.A(\count_cycle[19] ),
    .B(\count_cycle[20] ),
    .C(_06932_),
    .X(_06935_));
 sky130_fd_sc_hd__a21o_1 _27653_ (.A1(\count_cycle[19] ),
    .A2(_06932_),
    .B1(\count_cycle[20] ),
    .X(_06936_));
 sky130_fd_sc_hd__and3b_1 _27654_ (.A_N(_06935_),
    .B(_06916_),
    .C(_06936_),
    .X(_06937_));
 sky130_fd_sc_hd__clkbuf_1 _27655_ (.A(_06937_),
    .X(_00955_));
 sky130_fd_sc_hd__and4_1 _27656_ (.A(\count_cycle[19] ),
    .B(\count_cycle[20] ),
    .C(\count_cycle[21] ),
    .D(_06932_),
    .X(_06938_));
 sky130_fd_sc_hd__o21ai_1 _27657_ (.A1(\count_cycle[21] ),
    .A2(_06935_),
    .B1(_06926_),
    .Y(_06939_));
 sky130_fd_sc_hd__nor2_1 _27658_ (.A(_06938_),
    .B(_06939_),
    .Y(_00956_));
 sky130_fd_sc_hd__a21oi_1 _27659_ (.A1(\count_cycle[22] ),
    .A2(_06938_),
    .B1(_06907_),
    .Y(_06940_));
 sky130_fd_sc_hd__o21a_1 _27660_ (.A1(\count_cycle[22] ),
    .A2(_06938_),
    .B1(_06940_),
    .X(_00957_));
 sky130_fd_sc_hd__and3_1 _27661_ (.A(\count_cycle[22] ),
    .B(\count_cycle[23] ),
    .C(_06938_),
    .X(_06941_));
 sky130_fd_sc_hd__a21o_1 _27662_ (.A1(\count_cycle[22] ),
    .A2(_06938_),
    .B1(\count_cycle[23] ),
    .X(_06942_));
 sky130_fd_sc_hd__and3b_1 _27663_ (.A_N(_06941_),
    .B(_06916_),
    .C(_06942_),
    .X(_06943_));
 sky130_fd_sc_hd__clkbuf_1 _27664_ (.A(_06943_),
    .X(_00958_));
 sky130_fd_sc_hd__and4_2 _27665_ (.A(\count_cycle[22] ),
    .B(\count_cycle[23] ),
    .C(\count_cycle[24] ),
    .D(_06938_),
    .X(_06944_));
 sky130_fd_sc_hd__o21ai_1 _27666_ (.A1(\count_cycle[24] ),
    .A2(_06941_),
    .B1(_06926_),
    .Y(_06945_));
 sky130_fd_sc_hd__nor2_1 _27667_ (.A(_06944_),
    .B(_06945_),
    .Y(_00959_));
 sky130_fd_sc_hd__buf_2 _27668_ (.A(_08183_),
    .X(_06946_));
 sky130_fd_sc_hd__a21oi_1 _27669_ (.A1(\count_cycle[25] ),
    .A2(_06944_),
    .B1(_06946_),
    .Y(_06947_));
 sky130_fd_sc_hd__o21a_1 _27670_ (.A1(\count_cycle[25] ),
    .A2(_06944_),
    .B1(_06947_),
    .X(_00960_));
 sky130_fd_sc_hd__and3_1 _27671_ (.A(\count_cycle[25] ),
    .B(\count_cycle[26] ),
    .C(_06944_),
    .X(_06948_));
 sky130_fd_sc_hd__a21o_1 _27672_ (.A1(\count_cycle[25] ),
    .A2(_06944_),
    .B1(\count_cycle[26] ),
    .X(_06949_));
 sky130_fd_sc_hd__and3b_1 _27673_ (.A_N(_06948_),
    .B(_06916_),
    .C(_06949_),
    .X(_06950_));
 sky130_fd_sc_hd__clkbuf_1 _27674_ (.A(_06950_),
    .X(_00961_));
 sky130_fd_sc_hd__and4_2 _27675_ (.A(\count_cycle[25] ),
    .B(\count_cycle[26] ),
    .C(\count_cycle[27] ),
    .D(_06944_),
    .X(_06951_));
 sky130_fd_sc_hd__o21ai_1 _27676_ (.A1(\count_cycle[27] ),
    .A2(_06948_),
    .B1(_06926_),
    .Y(_06952_));
 sky130_fd_sc_hd__nor2_1 _27677_ (.A(_06951_),
    .B(_06952_),
    .Y(_00962_));
 sky130_fd_sc_hd__a21oi_1 _27678_ (.A1(\count_cycle[28] ),
    .A2(_06951_),
    .B1(_06946_),
    .Y(_06953_));
 sky130_fd_sc_hd__o21a_1 _27679_ (.A1(\count_cycle[28] ),
    .A2(_06951_),
    .B1(_06953_),
    .X(_00963_));
 sky130_fd_sc_hd__and3_1 _27680_ (.A(\count_cycle[28] ),
    .B(\count_cycle[29] ),
    .C(_06951_),
    .X(_06954_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27681_ (.A(_08505_),
    .X(_06955_));
 sky130_fd_sc_hd__a21o_1 _27682_ (.A1(\count_cycle[28] ),
    .A2(_06951_),
    .B1(\count_cycle[29] ),
    .X(_06956_));
 sky130_fd_sc_hd__and3b_1 _27683_ (.A_N(_06954_),
    .B(_06955_),
    .C(_06956_),
    .X(_06957_));
 sky130_fd_sc_hd__clkbuf_1 _27684_ (.A(_06957_),
    .X(_00964_));
 sky130_fd_sc_hd__and4_2 _27685_ (.A(\count_cycle[28] ),
    .B(\count_cycle[29] ),
    .C(\count_cycle[30] ),
    .D(_06951_),
    .X(_06958_));
 sky130_fd_sc_hd__o21ai_1 _27686_ (.A1(\count_cycle[30] ),
    .A2(_06954_),
    .B1(_06926_),
    .Y(_06959_));
 sky130_fd_sc_hd__nor2_1 _27687_ (.A(_06958_),
    .B(_06959_),
    .Y(_00965_));
 sky130_fd_sc_hd__a21oi_1 _27688_ (.A1(\count_cycle[31] ),
    .A2(_06958_),
    .B1(_06946_),
    .Y(_06960_));
 sky130_fd_sc_hd__o21a_1 _27689_ (.A1(\count_cycle[31] ),
    .A2(_06958_),
    .B1(_06960_),
    .X(_00966_));
 sky130_fd_sc_hd__and3_1 _27690_ (.A(\count_cycle[32] ),
    .B(\count_cycle[31] ),
    .C(_06958_),
    .X(_06961_));
 sky130_fd_sc_hd__a21o_1 _27691_ (.A1(\count_cycle[31] ),
    .A2(_06958_),
    .B1(\count_cycle[32] ),
    .X(_06962_));
 sky130_fd_sc_hd__and3b_1 _27692_ (.A_N(_06961_),
    .B(_06955_),
    .C(_06962_),
    .X(_06963_));
 sky130_fd_sc_hd__clkbuf_1 _27693_ (.A(_06963_),
    .X(_00967_));
 sky130_fd_sc_hd__and4_1 _27694_ (.A(\count_cycle[32] ),
    .B(\count_cycle[33] ),
    .C(\count_cycle[31] ),
    .D(_06958_),
    .X(_06964_));
 sky130_fd_sc_hd__clkbuf_2 _27695_ (.A(_06235_),
    .X(_06965_));
 sky130_fd_sc_hd__o21ai_1 _27696_ (.A1(\count_cycle[33] ),
    .A2(_06961_),
    .B1(_06965_),
    .Y(_06966_));
 sky130_fd_sc_hd__nor2_1 _27697_ (.A(_06964_),
    .B(_06966_),
    .Y(_00968_));
 sky130_fd_sc_hd__a21oi_1 _27698_ (.A1(\count_cycle[34] ),
    .A2(_06964_),
    .B1(_06946_),
    .Y(_06967_));
 sky130_fd_sc_hd__o21a_1 _27699_ (.A1(\count_cycle[34] ),
    .A2(_06964_),
    .B1(_06967_),
    .X(_00969_));
 sky130_fd_sc_hd__and3_1 _27700_ (.A(\count_cycle[34] ),
    .B(\count_cycle[35] ),
    .C(_06964_),
    .X(_06968_));
 sky130_fd_sc_hd__a21o_1 _27701_ (.A1(\count_cycle[34] ),
    .A2(_06964_),
    .B1(\count_cycle[35] ),
    .X(_06969_));
 sky130_fd_sc_hd__and3b_1 _27702_ (.A_N(_06968_),
    .B(_06955_),
    .C(_06969_),
    .X(_06970_));
 sky130_fd_sc_hd__clkbuf_1 _27703_ (.A(_06970_),
    .X(_00970_));
 sky130_fd_sc_hd__and4_2 _27704_ (.A(\count_cycle[34] ),
    .B(\count_cycle[35] ),
    .C(\count_cycle[36] ),
    .D(_06964_),
    .X(_06971_));
 sky130_fd_sc_hd__o21ai_1 _27705_ (.A1(\count_cycle[36] ),
    .A2(_06968_),
    .B1(_06965_),
    .Y(_06972_));
 sky130_fd_sc_hd__nor2_1 _27706_ (.A(_06971_),
    .B(_06972_),
    .Y(_00971_));
 sky130_fd_sc_hd__a21oi_1 _27707_ (.A1(\count_cycle[37] ),
    .A2(_06971_),
    .B1(_06946_),
    .Y(_06973_));
 sky130_fd_sc_hd__o21a_1 _27708_ (.A1(\count_cycle[37] ),
    .A2(_06971_),
    .B1(_06973_),
    .X(_00972_));
 sky130_fd_sc_hd__and3_1 _27709_ (.A(\count_cycle[37] ),
    .B(\count_cycle[38] ),
    .C(_06971_),
    .X(_06974_));
 sky130_fd_sc_hd__a21o_1 _27710_ (.A1(\count_cycle[37] ),
    .A2(_06971_),
    .B1(\count_cycle[38] ),
    .X(_06975_));
 sky130_fd_sc_hd__and3b_1 _27711_ (.A_N(_06974_),
    .B(_06955_),
    .C(_06975_),
    .X(_06976_));
 sky130_fd_sc_hd__clkbuf_1 _27712_ (.A(_06976_),
    .X(_00973_));
 sky130_fd_sc_hd__and4_1 _27713_ (.A(\count_cycle[37] ),
    .B(\count_cycle[38] ),
    .C(\count_cycle[39] ),
    .D(_06971_),
    .X(_06977_));
 sky130_fd_sc_hd__o21ai_1 _27714_ (.A1(\count_cycle[39] ),
    .A2(_06974_),
    .B1(_06965_),
    .Y(_06978_));
 sky130_fd_sc_hd__nor2_1 _27715_ (.A(_06977_),
    .B(_06978_),
    .Y(_00974_));
 sky130_fd_sc_hd__a21oi_1 _27716_ (.A1(\count_cycle[40] ),
    .A2(_06977_),
    .B1(_06946_),
    .Y(_06979_));
 sky130_fd_sc_hd__o21a_1 _27717_ (.A1(\count_cycle[40] ),
    .A2(_06977_),
    .B1(_06979_),
    .X(_00975_));
 sky130_fd_sc_hd__and3_1 _27718_ (.A(\count_cycle[40] ),
    .B(\count_cycle[41] ),
    .C(_06977_),
    .X(_06980_));
 sky130_fd_sc_hd__a21o_1 _27719_ (.A1(\count_cycle[40] ),
    .A2(_06977_),
    .B1(\count_cycle[41] ),
    .X(_06981_));
 sky130_fd_sc_hd__and3b_1 _27720_ (.A_N(_06980_),
    .B(_06955_),
    .C(_06981_),
    .X(_06982_));
 sky130_fd_sc_hd__clkbuf_1 _27721_ (.A(_06982_),
    .X(_00976_));
 sky130_fd_sc_hd__and2_1 _27722_ (.A(\count_cycle[42] ),
    .B(_06980_),
    .X(_06983_));
 sky130_fd_sc_hd__or2_1 _27723_ (.A(\count_cycle[42] ),
    .B(_06980_),
    .X(_06984_));
 sky130_fd_sc_hd__and3b_1 _27724_ (.A_N(_06983_),
    .B(_06955_),
    .C(_06984_),
    .X(_06985_));
 sky130_fd_sc_hd__clkbuf_1 _27725_ (.A(_06985_),
    .X(_00977_));
 sky130_fd_sc_hd__and3_1 _27726_ (.A(\count_cycle[42] ),
    .B(\count_cycle[43] ),
    .C(_06980_),
    .X(_06986_));
 sky130_fd_sc_hd__o21ai_1 _27727_ (.A1(\count_cycle[43] ),
    .A2(_06983_),
    .B1(_06965_),
    .Y(_06987_));
 sky130_fd_sc_hd__nor2_1 _27728_ (.A(_06986_),
    .B(_06987_),
    .Y(_00978_));
 sky130_fd_sc_hd__and3_1 _27729_ (.A(\count_cycle[43] ),
    .B(\count_cycle[44] ),
    .C(_06983_),
    .X(_06988_));
 sky130_fd_sc_hd__o21ai_1 _27730_ (.A1(\count_cycle[44] ),
    .A2(_06986_),
    .B1(_06965_),
    .Y(_06989_));
 sky130_fd_sc_hd__nor2_1 _27731_ (.A(_06988_),
    .B(_06989_),
    .Y(_00979_));
 sky130_fd_sc_hd__and2_1 _27732_ (.A(\count_cycle[45] ),
    .B(_06988_),
    .X(_06990_));
 sky130_fd_sc_hd__o21ai_1 _27733_ (.A1(\count_cycle[45] ),
    .A2(_06988_),
    .B1(_06965_),
    .Y(_06991_));
 sky130_fd_sc_hd__nor2_1 _27734_ (.A(_06990_),
    .B(_06991_),
    .Y(_00980_));
 sky130_fd_sc_hd__o21ai_1 _27735_ (.A1(\count_cycle[46] ),
    .A2(_06990_),
    .B1(_06180_),
    .Y(_06992_));
 sky130_fd_sc_hd__a21oi_1 _27736_ (.A1(\count_cycle[46] ),
    .A2(_06990_),
    .B1(_06992_),
    .Y(_00981_));
 sky130_fd_sc_hd__and3_1 _27737_ (.A(\count_cycle[46] ),
    .B(\count_cycle[47] ),
    .C(_06990_),
    .X(_06993_));
 sky130_fd_sc_hd__clkbuf_2 _27738_ (.A(_08505_),
    .X(_06994_));
 sky130_fd_sc_hd__a31o_1 _27739_ (.A1(\count_cycle[45] ),
    .A2(\count_cycle[46] ),
    .A3(_06988_),
    .B1(\count_cycle[47] ),
    .X(_06995_));
 sky130_fd_sc_hd__and3b_1 _27740_ (.A_N(_06993_),
    .B(_06994_),
    .C(_06995_),
    .X(_06996_));
 sky130_fd_sc_hd__clkbuf_1 _27741_ (.A(_06996_),
    .X(_00982_));
 sky130_fd_sc_hd__and2_1 _27742_ (.A(\count_cycle[48] ),
    .B(_06993_),
    .X(_06997_));
 sky130_fd_sc_hd__o21ai_1 _27743_ (.A1(\count_cycle[48] ),
    .A2(_06993_),
    .B1(_06328_),
    .Y(_06998_));
 sky130_fd_sc_hd__nor2_1 _27744_ (.A(_06997_),
    .B(_06998_),
    .Y(_00983_));
 sky130_fd_sc_hd__and3_1 _27745_ (.A(\count_cycle[48] ),
    .B(\count_cycle[49] ),
    .C(_06993_),
    .X(_06999_));
 sky130_fd_sc_hd__or2_1 _27746_ (.A(\count_cycle[49] ),
    .B(_06997_),
    .X(_07000_));
 sky130_fd_sc_hd__and3b_1 _27747_ (.A_N(_06999_),
    .B(_06994_),
    .C(_07000_),
    .X(_07001_));
 sky130_fd_sc_hd__clkbuf_1 _27748_ (.A(_07001_),
    .X(_00984_));
 sky130_fd_sc_hd__and2_1 _27749_ (.A(\count_cycle[50] ),
    .B(_06999_),
    .X(_07002_));
 sky130_fd_sc_hd__o21ai_1 _27750_ (.A1(\count_cycle[50] ),
    .A2(_06999_),
    .B1(_06328_),
    .Y(_07003_));
 sky130_fd_sc_hd__nor2_1 _27751_ (.A(_07002_),
    .B(_07003_),
    .Y(_00985_));
 sky130_fd_sc_hd__and3_1 _27752_ (.A(\count_cycle[50] ),
    .B(\count_cycle[51] ),
    .C(_06999_),
    .X(_07004_));
 sky130_fd_sc_hd__o21ai_1 _27753_ (.A1(\count_cycle[51] ),
    .A2(_07002_),
    .B1(_06328_),
    .Y(_07005_));
 sky130_fd_sc_hd__nor2_1 _27754_ (.A(_07004_),
    .B(_07005_),
    .Y(_00986_));
 sky130_fd_sc_hd__o21ai_1 _27755_ (.A1(\count_cycle[52] ),
    .A2(_07004_),
    .B1(_06180_),
    .Y(_07006_));
 sky130_fd_sc_hd__a21oi_1 _27756_ (.A1(\count_cycle[52] ),
    .A2(_07004_),
    .B1(_07006_),
    .Y(_00987_));
 sky130_fd_sc_hd__and3_1 _27757_ (.A(\count_cycle[52] ),
    .B(\count_cycle[53] ),
    .C(_07004_),
    .X(_07007_));
 sky130_fd_sc_hd__a21o_1 _27758_ (.A1(\count_cycle[52] ),
    .A2(_07004_),
    .B1(\count_cycle[53] ),
    .X(_07008_));
 sky130_fd_sc_hd__and3b_1 _27759_ (.A_N(_07007_),
    .B(_06994_),
    .C(_07008_),
    .X(_07009_));
 sky130_fd_sc_hd__clkbuf_1 _27760_ (.A(_07009_),
    .X(_00988_));
 sky130_fd_sc_hd__and2_1 _27761_ (.A(\count_cycle[54] ),
    .B(_07007_),
    .X(_07010_));
 sky130_fd_sc_hd__o21ai_1 _27762_ (.A1(\count_cycle[54] ),
    .A2(_07007_),
    .B1(_06328_),
    .Y(_07011_));
 sky130_fd_sc_hd__nor2_1 _27763_ (.A(_07010_),
    .B(_07011_),
    .Y(_00989_));
 sky130_fd_sc_hd__o21ai_1 _27764_ (.A1(\count_cycle[55] ),
    .A2(_07010_),
    .B1(_06180_),
    .Y(_07012_));
 sky130_fd_sc_hd__a21oi_1 _27765_ (.A1(\count_cycle[55] ),
    .A2(_07010_),
    .B1(_07012_),
    .Y(_00990_));
 sky130_fd_sc_hd__and3_1 _27766_ (.A(\count_cycle[55] ),
    .B(\count_cycle[56] ),
    .C(_07010_),
    .X(_07013_));
 sky130_fd_sc_hd__a31o_1 _27767_ (.A1(\count_cycle[54] ),
    .A2(\count_cycle[55] ),
    .A3(_07007_),
    .B1(\count_cycle[56] ),
    .X(_07014_));
 sky130_fd_sc_hd__and3b_1 _27768_ (.A_N(_07013_),
    .B(_06994_),
    .C(_07014_),
    .X(_07015_));
 sky130_fd_sc_hd__clkbuf_1 _27769_ (.A(_07015_),
    .X(_00991_));
 sky130_fd_sc_hd__and2_1 _27770_ (.A(\count_cycle[57] ),
    .B(_07013_),
    .X(_07016_));
 sky130_fd_sc_hd__or2_1 _27771_ (.A(\count_cycle[57] ),
    .B(_07013_),
    .X(_07017_));
 sky130_fd_sc_hd__and3b_1 _27772_ (.A_N(_07016_),
    .B(_06994_),
    .C(_07017_),
    .X(_07018_));
 sky130_fd_sc_hd__clkbuf_1 _27773_ (.A(_07018_),
    .X(_00992_));
 sky130_fd_sc_hd__a21oi_1 _27774_ (.A1(\count_cycle[58] ),
    .A2(_07016_),
    .B1(_08520_),
    .Y(_07019_));
 sky130_fd_sc_hd__o21a_1 _27775_ (.A1(\count_cycle[58] ),
    .A2(_07016_),
    .B1(_07019_),
    .X(_00993_));
 sky130_fd_sc_hd__and3_1 _27776_ (.A(\count_cycle[58] ),
    .B(\count_cycle[59] ),
    .C(_07016_),
    .X(_07020_));
 sky130_fd_sc_hd__a31o_1 _27777_ (.A1(\count_cycle[57] ),
    .A2(\count_cycle[58] ),
    .A3(_07013_),
    .B1(\count_cycle[59] ),
    .X(_07021_));
 sky130_fd_sc_hd__and3b_1 _27778_ (.A_N(_07020_),
    .B(_06994_),
    .C(_07021_),
    .X(_07022_));
 sky130_fd_sc_hd__clkbuf_1 _27779_ (.A(_07022_),
    .X(_00994_));
 sky130_fd_sc_hd__and2_1 _27780_ (.A(\count_cycle[60] ),
    .B(_07020_),
    .X(_07023_));
 sky130_fd_sc_hd__o21ai_1 _27781_ (.A1(\count_cycle[60] ),
    .A2(_07020_),
    .B1(_06328_),
    .Y(_07024_));
 sky130_fd_sc_hd__nor2_1 _27782_ (.A(_07023_),
    .B(_07024_),
    .Y(_00995_));
 sky130_fd_sc_hd__a21oi_1 _27783_ (.A1(\count_cycle[61] ),
    .A2(_07023_),
    .B1(_08520_),
    .Y(_07025_));
 sky130_fd_sc_hd__o21a_1 _27784_ (.A1(\count_cycle[61] ),
    .A2(_07023_),
    .B1(_07025_),
    .X(_00996_));
 sky130_fd_sc_hd__and3_1 _27785_ (.A(\count_cycle[61] ),
    .B(\count_cycle[62] ),
    .C(_07023_),
    .X(_07026_));
 sky130_fd_sc_hd__a31o_1 _27786_ (.A1(\count_cycle[60] ),
    .A2(\count_cycle[61] ),
    .A3(_07020_),
    .B1(\count_cycle[62] ),
    .X(_07027_));
 sky130_fd_sc_hd__and3b_1 _27787_ (.A_N(_07026_),
    .B(_08322_),
    .C(_07027_),
    .X(_07028_));
 sky130_fd_sc_hd__clkbuf_1 _27788_ (.A(_07028_),
    .X(_00997_));
 sky130_fd_sc_hd__o21ai_1 _27789_ (.A1(\count_cycle[63] ),
    .A2(_07026_),
    .B1(_06180_),
    .Y(_07029_));
 sky130_fd_sc_hd__a21oi_1 _27790_ (.A1(\count_cycle[63] ),
    .A2(_07026_),
    .B1(_07029_),
    .Y(_00998_));
 sky130_fd_sc_hd__clkbuf_2 _27791_ (.A(is_lui_auipc_jal),
    .X(_07030_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27792_ (.A(_07030_),
    .X(_07031_));
 sky130_fd_sc_hd__and2b_1 _27793_ (.A_N(instr_lui),
    .B(is_lui_auipc_jal),
    .X(_07032_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27794_ (.A(_07032_),
    .X(_07033_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27795_ (.A(_07033_),
    .X(_07034_));
 sky130_fd_sc_hd__a2bb2o_1 _27796_ (.A1_N(_07031_),
    .A2_N(_08635_),
    .B1(_07034_),
    .B2(_08667_),
    .X(_07035_));
 sky130_fd_sc_hd__xor2_1 _27797_ (.A(_08326_),
    .B(\decoded_imm[0] ),
    .X(_07036_));
 sky130_fd_sc_hd__mux2_1 _27798_ (.A0(_07035_),
    .A1(_07036_),
    .S(_08149_),
    .X(_07037_));
 sky130_fd_sc_hd__o21a_4 _27799_ (.A1(_08178_),
    .A2(_08148_),
    .B1(_08172_),
    .X(_07038_));
 sky130_fd_sc_hd__buf_2 _27800_ (.A(_07038_),
    .X(_07039_));
 sky130_fd_sc_hd__mux2_1 _27801_ (.A0(_10264_),
    .A1(_07037_),
    .S(_07039_),
    .X(_07040_));
 sky130_fd_sc_hd__clkbuf_1 _27802_ (.A(_07040_),
    .X(_00999_));
 sky130_fd_sc_hd__o21ai_4 _27803_ (.A1(_08945_),
    .A2(_08149_),
    .B1(_08172_),
    .Y(_07041_));
 sky130_fd_sc_hd__clkbuf_4 _27804_ (.A(_08149_),
    .X(_07042_));
 sky130_fd_sc_hd__clkbuf_2 _27805_ (.A(_07030_),
    .X(_07043_));
 sky130_fd_sc_hd__clkbuf_2 _27806_ (.A(_07033_),
    .X(_07044_));
 sky130_fd_sc_hd__a2bb2o_1 _27807_ (.A1_N(_07043_),
    .A2_N(_08744_),
    .B1(_07044_),
    .B2(_08184_),
    .X(_07045_));
 sky130_fd_sc_hd__xor2_1 _27808_ (.A(net278),
    .B(\decoded_imm[1] ),
    .X(_07046_));
 sky130_fd_sc_hd__and3_1 _27809_ (.A(_08326_),
    .B(_08668_),
    .C(_07046_),
    .X(_07047_));
 sky130_fd_sc_hd__a21oi_1 _27810_ (.A1(_10264_),
    .A2(_08668_),
    .B1(_07046_),
    .Y(_07048_));
 sky130_fd_sc_hd__buf_2 _27811_ (.A(_08148_),
    .X(_07049_));
 sky130_fd_sc_hd__o21ai_1 _27812_ (.A1(_07047_),
    .A2(_07048_),
    .B1(_07049_),
    .Y(_07050_));
 sky130_fd_sc_hd__o211a_1 _27813_ (.A1(_07042_),
    .A2(_07045_),
    .B1(_07050_),
    .C1(_07039_),
    .X(_07051_));
 sky130_fd_sc_hd__a21o_1 _27814_ (.A1(_10104_),
    .A2(_07041_),
    .B1(_07051_),
    .X(_01000_));
 sky130_fd_sc_hd__a2bb2o_1 _27815_ (.A1_N(_07043_),
    .A2_N(_08798_),
    .B1(_07044_),
    .B2(_05008_),
    .X(_07052_));
 sky130_fd_sc_hd__nand2_1 _27816_ (.A(net289),
    .B(\decoded_imm[2] ),
    .Y(_07053_));
 sky130_fd_sc_hd__or2_1 _27817_ (.A(net289),
    .B(\decoded_imm[2] ),
    .X(_07054_));
 sky130_fd_sc_hd__and2_1 _27818_ (.A(net278),
    .B(_08762_),
    .X(_07055_));
 sky130_fd_sc_hd__a31o_1 _27819_ (.A1(net267),
    .A2(\decoded_imm[0] ),
    .A3(_07046_),
    .B1(_07055_),
    .X(_07056_));
 sky130_fd_sc_hd__and3_1 _27820_ (.A(_07053_),
    .B(_07054_),
    .C(_07056_),
    .X(_07057_));
 sky130_fd_sc_hd__a21oi_1 _27821_ (.A1(_07053_),
    .A2(_07054_),
    .B1(_07056_),
    .Y(_07058_));
 sky130_fd_sc_hd__o21ai_1 _27822_ (.A1(_07057_),
    .A2(_07058_),
    .B1(_07049_),
    .Y(_07059_));
 sky130_fd_sc_hd__o211a_1 _27823_ (.A1(_07042_),
    .A2(_07052_),
    .B1(_07059_),
    .C1(_07039_),
    .X(_07060_));
 sky130_fd_sc_hd__a21o_1 _27824_ (.A1(_10311_),
    .A2(_07041_),
    .B1(_07060_),
    .X(_01001_));
 sky130_fd_sc_hd__buf_1 _27825_ (.A(_07030_),
    .X(_07061_));
 sky130_fd_sc_hd__buf_1 _27826_ (.A(_07033_),
    .X(_07062_));
 sky130_fd_sc_hd__a2bb2o_1 _27827_ (.A1_N(_07061_),
    .A2_N(_08865_),
    .B1(_07062_),
    .B2(_08874_),
    .X(_07063_));
 sky130_fd_sc_hd__nand2_1 _27828_ (.A(net292),
    .B(\decoded_imm[3] ),
    .Y(_07064_));
 sky130_fd_sc_hd__or2_1 _27829_ (.A(net292),
    .B(\decoded_imm[3] ),
    .X(_07065_));
 sky130_fd_sc_hd__nand2_1 _27830_ (.A(_07064_),
    .B(_07065_),
    .Y(_07066_));
 sky130_fd_sc_hd__a21bo_1 _27831_ (.A1(_07054_),
    .A2(_07056_),
    .B1_N(_07053_),
    .X(_07067_));
 sky130_fd_sc_hd__xnor2_1 _27832_ (.A(_07066_),
    .B(_07067_),
    .Y(_07068_));
 sky130_fd_sc_hd__mux2_1 _27833_ (.A0(_07063_),
    .A1(_07068_),
    .S(_08149_),
    .X(_07069_));
 sky130_fd_sc_hd__mux2_1 _27834_ (.A0(_10322_),
    .A1(_07069_),
    .S(_07039_),
    .X(_07070_));
 sky130_fd_sc_hd__clkbuf_1 _27835_ (.A(_07070_),
    .X(_01002_));
 sky130_fd_sc_hd__nor2_1 _27836_ (.A(_07043_),
    .B(_08934_),
    .Y(_07071_));
 sky130_fd_sc_hd__a211o_1 _27837_ (.A1(\reg_pc[4] ),
    .A2(_07044_),
    .B1(_07071_),
    .C1(_07042_),
    .X(_07072_));
 sky130_fd_sc_hd__nand2_1 _27838_ (.A(net293),
    .B(\decoded_imm[4] ),
    .Y(_07073_));
 sky130_fd_sc_hd__or2_1 _27839_ (.A(net293),
    .B(\decoded_imm[4] ),
    .X(_07074_));
 sky130_fd_sc_hd__nand2_1 _27840_ (.A(_07073_),
    .B(_07074_),
    .Y(_07075_));
 sky130_fd_sc_hd__a21bo_1 _27841_ (.A1(_07065_),
    .A2(_07067_),
    .B1_N(_07064_),
    .X(_07076_));
 sky130_fd_sc_hd__xor2_1 _27842_ (.A(_07075_),
    .B(_07076_),
    .X(_07077_));
 sky130_fd_sc_hd__a21oi_1 _27843_ (.A1(_07042_),
    .A2(_07077_),
    .B1(_07041_),
    .Y(_07078_));
 sky130_fd_sc_hd__a22o_1 _27844_ (.A1(_10331_),
    .A2(_07041_),
    .B1(_07072_),
    .B2(_07078_),
    .X(_01003_));
 sky130_fd_sc_hd__nor2_1 _27845_ (.A(net294),
    .B(\decoded_imm[5] ),
    .Y(_07079_));
 sky130_fd_sc_hd__and2_1 _27846_ (.A(net294),
    .B(\decoded_imm[5] ),
    .X(_07080_));
 sky130_vsdinv _27847_ (.A(_07073_),
    .Y(_07081_));
 sky130_fd_sc_hd__a21oi_1 _27848_ (.A1(_07074_),
    .A2(_07076_),
    .B1(_07081_),
    .Y(_07082_));
 sky130_fd_sc_hd__o21ai_1 _27849_ (.A1(_07079_),
    .A2(_07080_),
    .B1(_07082_),
    .Y(_07083_));
 sky130_fd_sc_hd__or3_1 _27850_ (.A(_07082_),
    .B(_07079_),
    .C(_07080_),
    .X(_07084_));
 sky130_fd_sc_hd__clkbuf_2 _27851_ (.A(_07032_),
    .X(_07085_));
 sky130_fd_sc_hd__o2bb2a_1 _27852_ (.A1_N(\reg_pc[5] ),
    .A2_N(_07085_),
    .B1(_08978_),
    .B2(_07030_),
    .X(_07086_));
 sky130_fd_sc_hd__nor2_1 _27853_ (.A(_08149_),
    .B(_07086_),
    .Y(_07087_));
 sky130_fd_sc_hd__a31o_1 _27854_ (.A1(_07049_),
    .A2(_07083_),
    .A3(_07084_),
    .B1(_07087_),
    .X(_07088_));
 sky130_fd_sc_hd__mux2_1 _27855_ (.A0(_10334_),
    .A1(_07088_),
    .S(_07039_),
    .X(_07089_));
 sky130_fd_sc_hd__clkbuf_1 _27856_ (.A(_07089_),
    .X(_01004_));
 sky130_fd_sc_hd__nand2_1 _27857_ (.A(net295),
    .B(\decoded_imm[6] ),
    .Y(_07090_));
 sky130_fd_sc_hd__or2_1 _27858_ (.A(net295),
    .B(\decoded_imm[6] ),
    .X(_07091_));
 sky130_fd_sc_hd__nand2_1 _27859_ (.A(_07090_),
    .B(_07091_),
    .Y(_07092_));
 sky130_fd_sc_hd__a211oi_2 _27860_ (.A1(_07074_),
    .A2(_07076_),
    .B1(_07080_),
    .C1(_07081_),
    .Y(_07093_));
 sky130_fd_sc_hd__nor2_1 _27861_ (.A(_07079_),
    .B(_07093_),
    .Y(_07094_));
 sky130_fd_sc_hd__xor2_1 _27862_ (.A(_07092_),
    .B(_07094_),
    .X(_07095_));
 sky130_fd_sc_hd__nand2_1 _27863_ (.A(_08997_),
    .B(_07044_),
    .Y(_07096_));
 sky130_fd_sc_hd__o211a_1 _27864_ (.A1(_07043_),
    .A2(_09033_),
    .B1(_07096_),
    .C1(_08526_),
    .X(_07097_));
 sky130_fd_sc_hd__a21oi_1 _27865_ (.A1(_07049_),
    .A2(_07095_),
    .B1(_07097_),
    .Y(_07098_));
 sky130_fd_sc_hd__mux2_1 _27866_ (.A0(_10337_),
    .A1(_07098_),
    .S(_07039_),
    .X(_07099_));
 sky130_fd_sc_hd__clkbuf_1 _27867_ (.A(_07099_),
    .X(_01005_));
 sky130_fd_sc_hd__nand2_1 _27868_ (.A(net296),
    .B(\decoded_imm[7] ),
    .Y(_07100_));
 sky130_fd_sc_hd__or2_1 _27869_ (.A(net296),
    .B(\decoded_imm[7] ),
    .X(_07101_));
 sky130_fd_sc_hd__nand2_1 _27870_ (.A(_07100_),
    .B(_07101_),
    .Y(_07102_));
 sky130_fd_sc_hd__o31ai_2 _27871_ (.A1(_07079_),
    .A2(_07092_),
    .A3(_07093_),
    .B1(_07090_),
    .Y(_07103_));
 sky130_fd_sc_hd__xnor2_1 _27872_ (.A(_07102_),
    .B(_07103_),
    .Y(_07104_));
 sky130_fd_sc_hd__a2bb2o_1 _27873_ (.A1_N(_07061_),
    .A2_N(_09093_),
    .B1(_07062_),
    .B2(\reg_pc[7] ),
    .X(_07105_));
 sky130_fd_sc_hd__buf_2 _27874_ (.A(_08291_),
    .X(_07106_));
 sky130_fd_sc_hd__mux2_1 _27875_ (.A0(_07104_),
    .A1(_07105_),
    .S(_07106_),
    .X(_07107_));
 sky130_fd_sc_hd__clkbuf_2 _27876_ (.A(_07038_),
    .X(_07108_));
 sky130_fd_sc_hd__mux2_1 _27877_ (.A0(_08461_),
    .A1(_07107_),
    .S(_07108_),
    .X(_07109_));
 sky130_fd_sc_hd__clkbuf_1 _27878_ (.A(_07109_),
    .X(_01006_));
 sky130_fd_sc_hd__nand2_1 _27879_ (.A(net297),
    .B(\decoded_imm[8] ),
    .Y(_07110_));
 sky130_fd_sc_hd__or2_1 _27880_ (.A(net297),
    .B(\decoded_imm[8] ),
    .X(_07111_));
 sky130_fd_sc_hd__nand2_1 _27881_ (.A(_07110_),
    .B(_07111_),
    .Y(_07112_));
 sky130_fd_sc_hd__a21boi_1 _27882_ (.A1(_07101_),
    .A2(_07103_),
    .B1_N(_07100_),
    .Y(_07113_));
 sky130_fd_sc_hd__xor2_1 _27883_ (.A(_07112_),
    .B(_07113_),
    .X(_07114_));
 sky130_fd_sc_hd__a2bb2o_1 _27884_ (.A1_N(_07061_),
    .A2_N(_09151_),
    .B1(_07062_),
    .B2(\reg_pc[8] ),
    .X(_07115_));
 sky130_fd_sc_hd__mux2_1 _27885_ (.A0(_07114_),
    .A1(_07115_),
    .S(_07106_),
    .X(_07116_));
 sky130_fd_sc_hd__mux2_1 _27886_ (.A0(_10344_),
    .A1(_07116_),
    .S(_07108_),
    .X(_07117_));
 sky130_fd_sc_hd__clkbuf_1 _27887_ (.A(_07117_),
    .X(_01007_));
 sky130_fd_sc_hd__o21a_1 _27888_ (.A1(_07112_),
    .A2(_07113_),
    .B1(_07110_),
    .X(_07118_));
 sky130_fd_sc_hd__nand2_1 _27889_ (.A(net298),
    .B(\decoded_imm[9] ),
    .Y(_07119_));
 sky130_vsdinv _27890_ (.A(_07119_),
    .Y(_07120_));
 sky130_fd_sc_hd__nor2_1 _27891_ (.A(net298),
    .B(\decoded_imm[9] ),
    .Y(_07121_));
 sky130_fd_sc_hd__nor2_1 _27892_ (.A(_07120_),
    .B(_07121_),
    .Y(_07122_));
 sky130_fd_sc_hd__xnor2_1 _27893_ (.A(_07118_),
    .B(_07122_),
    .Y(_07123_));
 sky130_fd_sc_hd__a2bb2o_1 _27894_ (.A1_N(_07061_),
    .A2_N(_09205_),
    .B1(_07062_),
    .B2(_09170_),
    .X(_07124_));
 sky130_fd_sc_hd__mux2_1 _27895_ (.A0(_07123_),
    .A1(_07124_),
    .S(_07106_),
    .X(_07125_));
 sky130_fd_sc_hd__mux2_1 _27896_ (.A0(_10157_),
    .A1(_07125_),
    .S(_07108_),
    .X(_07126_));
 sky130_fd_sc_hd__clkbuf_1 _27897_ (.A(_07126_),
    .X(_01008_));
 sky130_fd_sc_hd__or2_1 _27898_ (.A(net268),
    .B(\decoded_imm[10] ),
    .X(_07127_));
 sky130_fd_sc_hd__nand2_1 _27899_ (.A(net268),
    .B(_09219_),
    .Y(_07128_));
 sky130_fd_sc_hd__nand2_1 _27900_ (.A(_07127_),
    .B(_07128_),
    .Y(_07129_));
 sky130_fd_sc_hd__a211o_1 _27901_ (.A1(_07118_),
    .A2(_07119_),
    .B1(_07121_),
    .C1(_07129_),
    .X(_07130_));
 sky130_fd_sc_hd__a21o_1 _27902_ (.A1(_07118_),
    .A2(_07119_),
    .B1(_07121_),
    .X(_07131_));
 sky130_fd_sc_hd__nand2_1 _27903_ (.A(_07129_),
    .B(_07131_),
    .Y(_07132_));
 sky130_fd_sc_hd__and2_1 _27904_ (.A(_07130_),
    .B(_07132_),
    .X(_07133_));
 sky130_fd_sc_hd__a2bb2o_1 _27905_ (.A1_N(_07061_),
    .A2_N(_09245_),
    .B1(_07062_),
    .B2(_09218_),
    .X(_07134_));
 sky130_fd_sc_hd__mux2_1 _27906_ (.A0(_07133_),
    .A1(_07134_),
    .S(_07106_),
    .X(_07135_));
 sky130_fd_sc_hd__mux2_1 _27907_ (.A0(_10163_),
    .A1(_07135_),
    .S(_07108_),
    .X(_07136_));
 sky130_fd_sc_hd__clkbuf_1 _27908_ (.A(_07136_),
    .X(_01009_));
 sky130_fd_sc_hd__nor2_1 _27909_ (.A(net269),
    .B(\decoded_imm[11] ),
    .Y(_07137_));
 sky130_fd_sc_hd__nand2_1 _27910_ (.A(net269),
    .B(\decoded_imm[11] ),
    .Y(_07138_));
 sky130_fd_sc_hd__or2b_1 _27911_ (.A(_07137_),
    .B_N(_07138_),
    .X(_07139_));
 sky130_fd_sc_hd__a21oi_1 _27912_ (.A1(_07128_),
    .A2(_07130_),
    .B1(_07139_),
    .Y(_07140_));
 sky130_fd_sc_hd__a31o_1 _27913_ (.A1(_07128_),
    .A2(_07130_),
    .A3(_07139_),
    .B1(_08526_),
    .X(_07141_));
 sky130_fd_sc_hd__a2bb2o_1 _27914_ (.A1_N(_07031_),
    .A2_N(_09282_),
    .B1(_07034_),
    .B2(_09295_),
    .X(_07142_));
 sky130_fd_sc_hd__a2bb2o_1 _27915_ (.A1_N(_07140_),
    .A2_N(_07141_),
    .B1(_07142_),
    .B2(_08527_),
    .X(_07143_));
 sky130_fd_sc_hd__mux2_1 _27916_ (.A0(_08412_),
    .A1(_07143_),
    .S(_07108_),
    .X(_07144_));
 sky130_fd_sc_hd__clkbuf_1 _27917_ (.A(_07144_),
    .X(_01010_));
 sky130_fd_sc_hd__or2_1 _27918_ (.A(net270),
    .B(\decoded_imm[12] ),
    .X(_07145_));
 sky130_fd_sc_hd__nand2_1 _27919_ (.A(net270),
    .B(_09305_),
    .Y(_07146_));
 sky130_fd_sc_hd__nand2_1 _27920_ (.A(_07145_),
    .B(_07146_),
    .Y(_07147_));
 sky130_fd_sc_hd__a31oi_1 _27921_ (.A1(_07128_),
    .A2(_07130_),
    .A3(_07138_),
    .B1(_07137_),
    .Y(_07148_));
 sky130_fd_sc_hd__xnor2_1 _27922_ (.A(_07147_),
    .B(_07148_),
    .Y(_07149_));
 sky130_fd_sc_hd__a2bb2o_1 _27923_ (.A1_N(_07061_),
    .A2_N(_09332_),
    .B1(_07062_),
    .B2(_09347_),
    .X(_07150_));
 sky130_fd_sc_hd__buf_2 _27924_ (.A(_08291_),
    .X(_07151_));
 sky130_fd_sc_hd__mux2_1 _27925_ (.A0(_07149_),
    .A1(_07150_),
    .S(_07151_),
    .X(_07152_));
 sky130_fd_sc_hd__mux2_1 _27926_ (.A0(_10354_),
    .A1(_07152_),
    .S(_07108_),
    .X(_07153_));
 sky130_fd_sc_hd__clkbuf_1 _27927_ (.A(_07153_),
    .X(_01011_));
 sky130_fd_sc_hd__nor2_1 _27928_ (.A(net271),
    .B(\decoded_imm[13] ),
    .Y(_07154_));
 sky130_fd_sc_hd__nand2_1 _27929_ (.A(net271),
    .B(\decoded_imm[13] ),
    .Y(_07155_));
 sky130_fd_sc_hd__or2b_1 _27930_ (.A(_07154_),
    .B_N(_07155_),
    .X(_07156_));
 sky130_fd_sc_hd__or2b_1 _27931_ (.A(_07147_),
    .B_N(_07148_),
    .X(_07157_));
 sky130_fd_sc_hd__nand2_1 _27932_ (.A(_07146_),
    .B(_07157_),
    .Y(_07158_));
 sky130_fd_sc_hd__xnor2_1 _27933_ (.A(_07156_),
    .B(_07158_),
    .Y(_07159_));
 sky130_fd_sc_hd__buf_1 _27934_ (.A(is_lui_auipc_jal),
    .X(_07160_));
 sky130_fd_sc_hd__buf_1 _27935_ (.A(_07033_),
    .X(_07161_));
 sky130_fd_sc_hd__a2bb2o_1 _27936_ (.A1_N(_07160_),
    .A2_N(_09372_),
    .B1(_07161_),
    .B2(\reg_pc[13] ),
    .X(_07162_));
 sky130_fd_sc_hd__mux2_1 _27937_ (.A0(_07159_),
    .A1(_07162_),
    .S(_07151_),
    .X(_07163_));
 sky130_fd_sc_hd__clkbuf_2 _27938_ (.A(_07038_),
    .X(_07164_));
 sky130_fd_sc_hd__mux2_1 _27939_ (.A0(_10357_),
    .A1(_07163_),
    .S(_07164_),
    .X(_07165_));
 sky130_fd_sc_hd__clkbuf_1 _27940_ (.A(_07165_),
    .X(_01012_));
 sky130_fd_sc_hd__or2_1 _27941_ (.A(net272),
    .B(\decoded_imm[14] ),
    .X(_07166_));
 sky130_fd_sc_hd__nand2_1 _27942_ (.A(net272),
    .B(\decoded_imm[14] ),
    .Y(_07167_));
 sky130_fd_sc_hd__nand2_1 _27943_ (.A(_07166_),
    .B(_07167_),
    .Y(_07168_));
 sky130_fd_sc_hd__a311o_1 _27944_ (.A1(_07146_),
    .A2(_07157_),
    .A3(_07155_),
    .B1(_07168_),
    .C1(_07154_),
    .X(_07169_));
 sky130_fd_sc_hd__a31o_1 _27945_ (.A1(_07146_),
    .A2(_07157_),
    .A3(_07155_),
    .B1(_07154_),
    .X(_07170_));
 sky130_fd_sc_hd__nand2_1 _27946_ (.A(_07168_),
    .B(_07170_),
    .Y(_07171_));
 sky130_fd_sc_hd__nand2_1 _27947_ (.A(_07169_),
    .B(_07171_),
    .Y(_07172_));
 sky130_fd_sc_hd__nand2_1 _27948_ (.A(_09386_),
    .B(_07044_),
    .Y(_07173_));
 sky130_fd_sc_hd__o211a_1 _27949_ (.A1(_07043_),
    .A2(_09414_),
    .B1(_07173_),
    .C1(_08527_),
    .X(_07174_));
 sky130_fd_sc_hd__a211o_1 _27950_ (.A1(_07042_),
    .A2(_07172_),
    .B1(_07174_),
    .C1(_07041_),
    .X(_07175_));
 sky130_fd_sc_hd__a21bo_1 _27951_ (.A1(_10361_),
    .A2(_07041_),
    .B1_N(_07175_),
    .X(_01013_));
 sky130_fd_sc_hd__nor2_1 _27952_ (.A(net273),
    .B(\decoded_imm[15] ),
    .Y(_07176_));
 sky130_fd_sc_hd__nand2_1 _27953_ (.A(net273),
    .B(\decoded_imm[15] ),
    .Y(_07177_));
 sky130_fd_sc_hd__or2b_1 _27954_ (.A(_07176_),
    .B_N(_07177_),
    .X(_07178_));
 sky130_fd_sc_hd__a21oi_1 _27955_ (.A1(_07167_),
    .A2(_07169_),
    .B1(_07178_),
    .Y(_07179_));
 sky130_fd_sc_hd__a31o_1 _27956_ (.A1(_07167_),
    .A2(_07169_),
    .A3(_07178_),
    .B1(_08526_),
    .X(_07180_));
 sky130_fd_sc_hd__a2bb2o_1 _27957_ (.A1_N(_07031_),
    .A2_N(_09453_),
    .B1(_07034_),
    .B2(\reg_pc[15] ),
    .X(_07181_));
 sky130_fd_sc_hd__a2bb2o_1 _27958_ (.A1_N(_07179_),
    .A2_N(_07180_),
    .B1(_07181_),
    .B2(_08527_),
    .X(_07182_));
 sky130_fd_sc_hd__mux2_1 _27959_ (.A0(_10187_),
    .A1(_07182_),
    .S(_07164_),
    .X(_07183_));
 sky130_fd_sc_hd__clkbuf_1 _27960_ (.A(_07183_),
    .X(_01014_));
 sky130_fd_sc_hd__or2_1 _27961_ (.A(net274),
    .B(\decoded_imm[16] ),
    .X(_07184_));
 sky130_fd_sc_hd__nand2_1 _27962_ (.A(net274),
    .B(\decoded_imm[16] ),
    .Y(_07185_));
 sky130_fd_sc_hd__nand2_1 _27963_ (.A(_07184_),
    .B(_07185_),
    .Y(_07186_));
 sky130_fd_sc_hd__a311o_1 _27964_ (.A1(_07167_),
    .A2(_07169_),
    .A3(_07177_),
    .B1(_07186_),
    .C1(_07176_),
    .X(_07187_));
 sky130_fd_sc_hd__a31o_1 _27965_ (.A1(_07167_),
    .A2(_07169_),
    .A3(_07177_),
    .B1(_07176_),
    .X(_07188_));
 sky130_fd_sc_hd__nand2_1 _27966_ (.A(_07186_),
    .B(_07188_),
    .Y(_07189_));
 sky130_fd_sc_hd__and2_1 _27967_ (.A(_07187_),
    .B(_07189_),
    .X(_07190_));
 sky130_fd_sc_hd__a2bb2o_1 _27968_ (.A1_N(_07160_),
    .A2_N(_09507_),
    .B1(_07161_),
    .B2(_09468_),
    .X(_07191_));
 sky130_fd_sc_hd__mux2_1 _27969_ (.A0(_07190_),
    .A1(_07191_),
    .S(_07151_),
    .X(_07192_));
 sky130_fd_sc_hd__mux2_1 _27970_ (.A0(_10367_),
    .A1(_07192_),
    .S(_07164_),
    .X(_07193_));
 sky130_fd_sc_hd__clkbuf_1 _27971_ (.A(_07193_),
    .X(_01015_));
 sky130_fd_sc_hd__nor2_1 _27972_ (.A(net275),
    .B(\decoded_imm[17] ),
    .Y(_07194_));
 sky130_fd_sc_hd__nand2_1 _27973_ (.A(net275),
    .B(\decoded_imm[17] ),
    .Y(_07195_));
 sky130_fd_sc_hd__or2b_1 _27974_ (.A(_07194_),
    .B_N(_07195_),
    .X(_07196_));
 sky130_fd_sc_hd__a21oi_1 _27975_ (.A1(_07185_),
    .A2(_07187_),
    .B1(_07196_),
    .Y(_07197_));
 sky130_fd_sc_hd__a31o_1 _27976_ (.A1(_07185_),
    .A2(_07187_),
    .A3(_07196_),
    .B1(_08526_),
    .X(_07198_));
 sky130_fd_sc_hd__a2bb2o_1 _27977_ (.A1_N(_07031_),
    .A2_N(_09545_),
    .B1(_07034_),
    .B2(\reg_pc[17] ),
    .X(_07199_));
 sky130_fd_sc_hd__a2bb2o_1 _27978_ (.A1_N(_07197_),
    .A2_N(_07198_),
    .B1(_07199_),
    .B2(_08527_),
    .X(_07200_));
 sky130_fd_sc_hd__mux2_1 _27979_ (.A0(_10197_),
    .A1(_07200_),
    .S(_07164_),
    .X(_07201_));
 sky130_fd_sc_hd__clkbuf_1 _27980_ (.A(_07201_),
    .X(_01016_));
 sky130_fd_sc_hd__or2_1 _27981_ (.A(net276),
    .B(\decoded_imm[18] ),
    .X(_07202_));
 sky130_fd_sc_hd__nand2_1 _27982_ (.A(net276),
    .B(\decoded_imm[18] ),
    .Y(_07203_));
 sky130_fd_sc_hd__nand2_1 _27983_ (.A(_07202_),
    .B(_07203_),
    .Y(_07204_));
 sky130_fd_sc_hd__a311o_1 _27984_ (.A1(_07185_),
    .A2(_07187_),
    .A3(_07195_),
    .B1(_07204_),
    .C1(_07194_),
    .X(_07205_));
 sky130_fd_sc_hd__a31o_1 _27985_ (.A1(_07185_),
    .A2(_07187_),
    .A3(_07195_),
    .B1(_07194_),
    .X(_07206_));
 sky130_fd_sc_hd__nand2_1 _27986_ (.A(_07204_),
    .B(_07206_),
    .Y(_07207_));
 sky130_fd_sc_hd__and2_1 _27987_ (.A(_07205_),
    .B(_07207_),
    .X(_07208_));
 sky130_fd_sc_hd__a2bb2o_1 _27988_ (.A1_N(_07160_),
    .A2_N(_09589_),
    .B1(_07161_),
    .B2(_05150_),
    .X(_07209_));
 sky130_fd_sc_hd__mux2_1 _27989_ (.A0(_07208_),
    .A1(_07209_),
    .S(_07151_),
    .X(_07210_));
 sky130_fd_sc_hd__mux2_1 _27990_ (.A0(_10372_),
    .A1(_07210_),
    .S(_07164_),
    .X(_07211_));
 sky130_fd_sc_hd__clkbuf_1 _27991_ (.A(_07211_),
    .X(_01017_));
 sky130_fd_sc_hd__nor2_1 _27992_ (.A(net277),
    .B(\decoded_imm[19] ),
    .Y(_07212_));
 sky130_fd_sc_hd__nand2_1 _27993_ (.A(net277),
    .B(\decoded_imm[19] ),
    .Y(_07213_));
 sky130_fd_sc_hd__or2b_1 _27994_ (.A(_07212_),
    .B_N(_07213_),
    .X(_07214_));
 sky130_fd_sc_hd__a21oi_1 _27995_ (.A1(_07203_),
    .A2(_07205_),
    .B1(_07214_),
    .Y(_07215_));
 sky130_fd_sc_hd__a31o_1 _27996_ (.A1(_07203_),
    .A2(_07205_),
    .A3(_07214_),
    .B1(_08291_),
    .X(_07216_));
 sky130_fd_sc_hd__a2bb2o_1 _27997_ (.A1_N(_07031_),
    .A2_N(_09626_),
    .B1(_07034_),
    .B2(\reg_pc[19] ),
    .X(_07217_));
 sky130_fd_sc_hd__a2bb2o_1 _27998_ (.A1_N(_07215_),
    .A2_N(_07216_),
    .B1(_07217_),
    .B2(_07106_),
    .X(_07218_));
 sky130_fd_sc_hd__mux2_1 _27999_ (.A0(_10206_),
    .A1(_07218_),
    .S(_07164_),
    .X(_07219_));
 sky130_fd_sc_hd__clkbuf_1 _28000_ (.A(_07219_),
    .X(_01018_));
 sky130_fd_sc_hd__or2_1 _28001_ (.A(net279),
    .B(\decoded_imm[20] ),
    .X(_07220_));
 sky130_fd_sc_hd__nand2_1 _28002_ (.A(net279),
    .B(\decoded_imm[20] ),
    .Y(_07221_));
 sky130_fd_sc_hd__nand2_1 _28003_ (.A(_07220_),
    .B(_07221_),
    .Y(_07222_));
 sky130_fd_sc_hd__a31o_1 _28004_ (.A1(_07203_),
    .A2(_07205_),
    .A3(_07213_),
    .B1(_07212_),
    .X(_07223_));
 sky130_fd_sc_hd__or2_1 _28005_ (.A(_07222_),
    .B(_07223_),
    .X(_07224_));
 sky130_fd_sc_hd__nand2_1 _28006_ (.A(_07222_),
    .B(_07223_),
    .Y(_07225_));
 sky130_fd_sc_hd__and2_1 _28007_ (.A(_07224_),
    .B(_07225_),
    .X(_07226_));
 sky130_fd_sc_hd__a2bb2o_1 _28008_ (.A1_N(_07160_),
    .A2_N(_09667_),
    .B1(_07161_),
    .B2(_09634_),
    .X(_07227_));
 sky130_fd_sc_hd__mux2_1 _28009_ (.A0(_07226_),
    .A1(_07227_),
    .S(_07151_),
    .X(_07228_));
 sky130_fd_sc_hd__clkbuf_2 _28010_ (.A(_07038_),
    .X(_07229_));
 sky130_fd_sc_hd__mux2_1 _28011_ (.A0(_10378_),
    .A1(_07228_),
    .S(_07229_),
    .X(_07230_));
 sky130_fd_sc_hd__clkbuf_1 _28012_ (.A(_07230_),
    .X(_01019_));
 sky130_fd_sc_hd__nor2_1 _28013_ (.A(net280),
    .B(\decoded_imm[21] ),
    .Y(_07231_));
 sky130_fd_sc_hd__nand2_1 _28014_ (.A(net280),
    .B(\decoded_imm[21] ),
    .Y(_07232_));
 sky130_fd_sc_hd__or2b_1 _28015_ (.A(_07231_),
    .B_N(_07232_),
    .X(_07233_));
 sky130_fd_sc_hd__a21oi_1 _28016_ (.A1(_07221_),
    .A2(_07224_),
    .B1(_07233_),
    .Y(_07234_));
 sky130_fd_sc_hd__a31o_1 _28017_ (.A1(_07221_),
    .A2(_07224_),
    .A3(_07233_),
    .B1(_08291_),
    .X(_07235_));
 sky130_fd_sc_hd__a2bb2o_1 _28018_ (.A1_N(_07031_),
    .A2_N(_09704_),
    .B1(_07034_),
    .B2(\reg_pc[21] ),
    .X(_07236_));
 sky130_fd_sc_hd__a2bb2o_1 _28019_ (.A1_N(_07234_),
    .A2_N(_07235_),
    .B1(_07236_),
    .B2(_07106_),
    .X(_07237_));
 sky130_fd_sc_hd__mux2_1 _28020_ (.A0(_10214_),
    .A1(_07237_),
    .S(_07229_),
    .X(_07238_));
 sky130_fd_sc_hd__clkbuf_1 _28021_ (.A(_07238_),
    .X(_01020_));
 sky130_fd_sc_hd__or2_1 _28022_ (.A(net281),
    .B(\decoded_imm[22] ),
    .X(_07239_));
 sky130_fd_sc_hd__nand2_1 _28023_ (.A(net281),
    .B(\decoded_imm[22] ),
    .Y(_07240_));
 sky130_fd_sc_hd__nand2_1 _28024_ (.A(_07239_),
    .B(_07240_),
    .Y(_07241_));
 sky130_fd_sc_hd__a31o_1 _28025_ (.A1(_07221_),
    .A2(_07224_),
    .A3(_07232_),
    .B1(_07231_),
    .X(_07242_));
 sky130_fd_sc_hd__xor2_1 _28026_ (.A(_07241_),
    .B(_07242_),
    .X(_07243_));
 sky130_fd_sc_hd__a2bb2o_1 _28027_ (.A1_N(_07160_),
    .A2_N(_09744_),
    .B1(_07161_),
    .B2(_09712_),
    .X(_07244_));
 sky130_fd_sc_hd__mux2_1 _28028_ (.A0(_07243_),
    .A1(_07244_),
    .S(_07151_),
    .X(_07245_));
 sky130_fd_sc_hd__mux2_1 _28029_ (.A0(_10384_),
    .A1(_07245_),
    .S(_07229_),
    .X(_07246_));
 sky130_fd_sc_hd__clkbuf_1 _28030_ (.A(_07246_),
    .X(_01021_));
 sky130_fd_sc_hd__or2_1 _28031_ (.A(net282),
    .B(\decoded_imm[23] ),
    .X(_07247_));
 sky130_fd_sc_hd__nand2_1 _28032_ (.A(_10223_),
    .B(_09751_),
    .Y(_07248_));
 sky130_fd_sc_hd__nand2_1 _28033_ (.A(_07247_),
    .B(_07248_),
    .Y(_07249_));
 sky130_fd_sc_hd__o21a_1 _28034_ (.A1(_07241_),
    .A2(_07242_),
    .B1(_07240_),
    .X(_07250_));
 sky130_fd_sc_hd__or2_1 _28035_ (.A(_07249_),
    .B(_07250_),
    .X(_07251_));
 sky130_fd_sc_hd__a21oi_1 _28036_ (.A1(_07249_),
    .A2(_07250_),
    .B1(_08526_),
    .Y(_07252_));
 sky130_fd_sc_hd__a2bb2o_1 _28037_ (.A1_N(_07043_),
    .A2_N(_09781_),
    .B1(_07044_),
    .B2(_09750_),
    .X(_07253_));
 sky130_fd_sc_hd__a22o_1 _28038_ (.A1(_07251_),
    .A2(_07252_),
    .B1(_07253_),
    .B2(_08527_),
    .X(_07254_));
 sky130_fd_sc_hd__mux2_1 _28039_ (.A0(_10224_),
    .A1(_07254_),
    .S(_07229_),
    .X(_07255_));
 sky130_fd_sc_hd__clkbuf_1 _28040_ (.A(_07255_),
    .X(_01022_));
 sky130_fd_sc_hd__and2_1 _28041_ (.A(net283),
    .B(\decoded_imm[24] ),
    .X(_07256_));
 sky130_fd_sc_hd__or2_1 _28042_ (.A(net283),
    .B(\decoded_imm[24] ),
    .X(_07257_));
 sky130_fd_sc_hd__or2b_1 _28043_ (.A(_07256_),
    .B_N(_07257_),
    .X(_07258_));
 sky130_fd_sc_hd__a21boi_1 _28044_ (.A1(_07248_),
    .A2(_07250_),
    .B1_N(_07247_),
    .Y(_07259_));
 sky130_fd_sc_hd__xnor2_1 _28045_ (.A(_07258_),
    .B(_07259_),
    .Y(_07260_));
 sky130_fd_sc_hd__a2bb2o_1 _28046_ (.A1_N(_07160_),
    .A2_N(_09821_),
    .B1(_07161_),
    .B2(_09788_),
    .X(_07261_));
 sky130_fd_sc_hd__clkbuf_2 _28047_ (.A(_08291_),
    .X(_07262_));
 sky130_fd_sc_hd__mux2_1 _28048_ (.A0(_07260_),
    .A1(_07261_),
    .S(_07262_),
    .X(_07263_));
 sky130_fd_sc_hd__mux2_1 _28049_ (.A0(_10389_),
    .A1(_07263_),
    .S(_07229_),
    .X(_07264_));
 sky130_fd_sc_hd__clkbuf_1 _28050_ (.A(_07264_),
    .X(_01023_));
 sky130_fd_sc_hd__a21o_1 _28051_ (.A1(_07257_),
    .A2(_07259_),
    .B1(_07256_),
    .X(_07265_));
 sky130_fd_sc_hd__or2_1 _28052_ (.A(net284),
    .B(\decoded_imm[25] ),
    .X(_07266_));
 sky130_fd_sc_hd__nand2_1 _28053_ (.A(_10232_),
    .B(\decoded_imm[25] ),
    .Y(_07267_));
 sky130_fd_sc_hd__nand2_1 _28054_ (.A(_07266_),
    .B(_07267_),
    .Y(_07268_));
 sky130_fd_sc_hd__xnor2_1 _28055_ (.A(_07265_),
    .B(_07268_),
    .Y(_07269_));
 sky130_fd_sc_hd__a2bb2o_1 _28056_ (.A1_N(_08496_),
    .A2_N(_09855_),
    .B1(_07085_),
    .B2(\reg_pc[25] ),
    .X(_07270_));
 sky130_fd_sc_hd__mux2_1 _28057_ (.A0(_07269_),
    .A1(_07270_),
    .S(_07262_),
    .X(_07271_));
 sky130_fd_sc_hd__mux2_1 _28058_ (.A0(_10392_),
    .A1(_07271_),
    .S(_07229_),
    .X(_07272_));
 sky130_fd_sc_hd__clkbuf_1 _28059_ (.A(_07272_),
    .X(_01024_));
 sky130_fd_sc_hd__nand2_1 _28060_ (.A(_10396_),
    .B(\decoded_imm[26] ),
    .Y(_07273_));
 sky130_fd_sc_hd__or2_1 _28061_ (.A(_10396_),
    .B(\decoded_imm[26] ),
    .X(_07274_));
 sky130_fd_sc_hd__nand2_1 _28062_ (.A(_07273_),
    .B(_07274_),
    .Y(_07275_));
 sky130_fd_sc_hd__a21boi_1 _28063_ (.A1(_07265_),
    .A2(_07266_),
    .B1_N(_07267_),
    .Y(_07276_));
 sky130_fd_sc_hd__xor2_1 _28064_ (.A(_07275_),
    .B(_07276_),
    .X(_07277_));
 sky130_fd_sc_hd__a2bb2o_1 _28065_ (.A1_N(_08496_),
    .A2_N(_09888_),
    .B1(_07085_),
    .B2(_09894_),
    .X(_07278_));
 sky130_fd_sc_hd__mux2_1 _28066_ (.A0(_07277_),
    .A1(_07278_),
    .S(_07262_),
    .X(_07279_));
 sky130_fd_sc_hd__buf_2 _28067_ (.A(_07038_),
    .X(_07280_));
 sky130_fd_sc_hd__mux2_1 _28068_ (.A0(_10397_),
    .A1(_07279_),
    .S(_07280_),
    .X(_07281_));
 sky130_fd_sc_hd__clkbuf_1 _28069_ (.A(_07281_),
    .X(_01025_));
 sky130_fd_sc_hd__o21a_1 _28070_ (.A1(_07275_),
    .A2(_07276_),
    .B1(_07273_),
    .X(_07282_));
 sky130_fd_sc_hd__nor2_1 _28071_ (.A(net286),
    .B(\decoded_imm[27] ),
    .Y(_07283_));
 sky130_fd_sc_hd__and2_1 _28072_ (.A(net286),
    .B(\decoded_imm[27] ),
    .X(_07284_));
 sky130_fd_sc_hd__or3_1 _28073_ (.A(_07282_),
    .B(_07283_),
    .C(_07284_),
    .X(_07285_));
 sky130_fd_sc_hd__o21ai_1 _28074_ (.A1(_07283_),
    .A2(_07284_),
    .B1(_07282_),
    .Y(_07286_));
 sky130_fd_sc_hd__o2bb2a_1 _28075_ (.A1_N(_09902_),
    .A2_N(_07033_),
    .B1(_09929_),
    .B2(_07030_),
    .X(_07287_));
 sky130_fd_sc_hd__nor2_1 _28076_ (.A(_08148_),
    .B(_07287_),
    .Y(_07288_));
 sky130_fd_sc_hd__a31o_1 _28077_ (.A1(_07049_),
    .A2(_07285_),
    .A3(_07286_),
    .B1(_07288_),
    .X(_07289_));
 sky130_fd_sc_hd__mux2_1 _28078_ (.A0(_10241_),
    .A1(_07289_),
    .S(_07280_),
    .X(_07290_));
 sky130_fd_sc_hd__clkbuf_1 _28079_ (.A(_07290_),
    .X(_01026_));
 sky130_fd_sc_hd__and2_1 _28080_ (.A(net287),
    .B(\decoded_imm[28] ),
    .X(_07291_));
 sky130_fd_sc_hd__or2_1 _28081_ (.A(net287),
    .B(\decoded_imm[28] ),
    .X(_07292_));
 sky130_fd_sc_hd__or2b_1 _28082_ (.A(_07291_),
    .B_N(_07292_),
    .X(_07293_));
 sky130_fd_sc_hd__o21bai_1 _28083_ (.A1(_07282_),
    .A2(_07283_),
    .B1_N(_07284_),
    .Y(_07294_));
 sky130_fd_sc_hd__xnor2_1 _28084_ (.A(_07293_),
    .B(_07294_),
    .Y(_07295_));
 sky130_fd_sc_hd__a2bb2o_1 _28085_ (.A1_N(_08496_),
    .A2_N(_09966_),
    .B1(_07085_),
    .B2(\reg_pc[28] ),
    .X(_07296_));
 sky130_fd_sc_hd__mux2_1 _28086_ (.A0(_07295_),
    .A1(_07296_),
    .S(_07262_),
    .X(_07297_));
 sky130_fd_sc_hd__mux2_1 _28087_ (.A0(_10246_),
    .A1(_07297_),
    .S(_07280_),
    .X(_07298_));
 sky130_fd_sc_hd__clkbuf_1 _28088_ (.A(_07298_),
    .X(_01027_));
 sky130_fd_sc_hd__a21oi_1 _28089_ (.A1(_07292_),
    .A2(_07294_),
    .B1(_07291_),
    .Y(_07299_));
 sky130_fd_sc_hd__nor2_1 _28090_ (.A(net288),
    .B(\decoded_imm[29] ),
    .Y(_07300_));
 sky130_fd_sc_hd__and2_1 _28091_ (.A(net288),
    .B(\decoded_imm[29] ),
    .X(_07301_));
 sky130_fd_sc_hd__or3_1 _28092_ (.A(_07299_),
    .B(_07300_),
    .C(_07301_),
    .X(_07302_));
 sky130_fd_sc_hd__o21ai_1 _28093_ (.A1(_07300_),
    .A2(_07301_),
    .B1(_07299_),
    .Y(_07303_));
 sky130_fd_sc_hd__o2bb2a_1 _28094_ (.A1_N(_09975_),
    .A2_N(_07033_),
    .B1(_10003_),
    .B2(_07030_),
    .X(_07304_));
 sky130_fd_sc_hd__nor2_1 _28095_ (.A(_08148_),
    .B(_07304_),
    .Y(_07305_));
 sky130_fd_sc_hd__a31o_1 _28096_ (.A1(_07049_),
    .A2(_07302_),
    .A3(_07303_),
    .B1(_07305_),
    .X(_07306_));
 sky130_fd_sc_hd__mux2_1 _28097_ (.A0(_10250_),
    .A1(_07306_),
    .S(_07280_),
    .X(_07307_));
 sky130_fd_sc_hd__clkbuf_1 _28098_ (.A(_07307_),
    .X(_01028_));
 sky130_fd_sc_hd__nand2_1 _28099_ (.A(_10254_),
    .B(\decoded_imm[30] ),
    .Y(_07308_));
 sky130_fd_sc_hd__or2_1 _28100_ (.A(net290),
    .B(\decoded_imm[30] ),
    .X(_07309_));
 sky130_fd_sc_hd__nand2_1 _28101_ (.A(_07308_),
    .B(_07309_),
    .Y(_07310_));
 sky130_fd_sc_hd__o21ba_1 _28102_ (.A1(_07299_),
    .A2(_07300_),
    .B1_N(_07301_),
    .X(_07311_));
 sky130_fd_sc_hd__xor2_1 _28103_ (.A(_07310_),
    .B(_07311_),
    .X(_07312_));
 sky130_fd_sc_hd__a2bb2o_1 _28104_ (.A1_N(_08496_),
    .A2_N(_10040_),
    .B1(_07085_),
    .B2(\reg_pc[30] ),
    .X(_07313_));
 sky130_fd_sc_hd__mux2_1 _28105_ (.A0(_07312_),
    .A1(_07313_),
    .S(_07262_),
    .X(_07314_));
 sky130_fd_sc_hd__mux2_1 _28106_ (.A0(_10255_),
    .A1(_07314_),
    .S(_07280_),
    .X(_07315_));
 sky130_fd_sc_hd__clkbuf_1 _28107_ (.A(_07315_),
    .X(_01029_));
 sky130_fd_sc_hd__o21ai_1 _28108_ (.A1(_07310_),
    .A2(_07311_),
    .B1(_07308_),
    .Y(_07316_));
 sky130_fd_sc_hd__xnor2_1 _28109_ (.A(_08393_),
    .B(\decoded_imm[31] ),
    .Y(_07317_));
 sky130_fd_sc_hd__xnor2_1 _28110_ (.A(_07316_),
    .B(_07317_),
    .Y(_07318_));
 sky130_fd_sc_hd__a2bb2o_1 _28111_ (.A1_N(_08496_),
    .A2_N(_10077_),
    .B1(_07085_),
    .B2(\reg_pc[31] ),
    .X(_07319_));
 sky130_fd_sc_hd__mux2_1 _28112_ (.A0(_07318_),
    .A1(_07319_),
    .S(_07262_),
    .X(_07320_));
 sky130_fd_sc_hd__mux2_1 _28113_ (.A0(_10259_),
    .A1(_07320_),
    .S(_07280_),
    .X(_07321_));
 sky130_fd_sc_hd__clkbuf_1 _28114_ (.A(_07321_),
    .X(_01030_));
 sky130_fd_sc_hd__or3_1 _28115_ (.A(_08186_),
    .B(_06117_),
    .C(_08280_),
    .X(_07322_));
 sky130_fd_sc_hd__o211a_1 _28116_ (.A1(irq_delay),
    .A2(_06182_),
    .B1(_07322_),
    .C1(_06175_),
    .X(_01031_));
 sky130_vsdinv _28117_ (.A(_04972_),
    .Y(_07323_));
 sky130_fd_sc_hd__nand2_1 _28118_ (.A(_07323_),
    .B(_08232_),
    .Y(_07324_));
 sky130_fd_sc_hd__nand2_1 _28119_ (.A(_06119_),
    .B(_07324_),
    .Y(_07325_));
 sky130_fd_sc_hd__a31o_1 _28120_ (.A1(_06118_),
    .A2(_06119_),
    .A3(_07324_),
    .B1(_08186_),
    .X(_07326_));
 sky130_fd_sc_hd__clkbuf_2 _28121_ (.A(_06179_),
    .X(_07327_));
 sky130_fd_sc_hd__buf_2 _28122_ (.A(_07327_),
    .X(_07328_));
 sky130_fd_sc_hd__o211a_1 _28123_ (.A1(_06126_),
    .A2(_07325_),
    .B1(_07326_),
    .C1(_07328_),
    .X(_01032_));
 sky130_fd_sc_hd__nand2_1 _28124_ (.A(_08179_),
    .B(_08638_),
    .Y(_07329_));
 sky130_fd_sc_hd__clkbuf_2 _28125_ (.A(_07329_),
    .X(_07330_));
 sky130_fd_sc_hd__clkbuf_2 _28126_ (.A(_07330_),
    .X(_07331_));
 sky130_fd_sc_hd__clkbuf_2 _28127_ (.A(_07329_),
    .X(_07332_));
 sky130_fd_sc_hd__nor2_1 _28128_ (.A(_08635_),
    .B(_07332_),
    .Y(_07333_));
 sky130_fd_sc_hd__clkbuf_2 _28129_ (.A(_08183_),
    .X(_07334_));
 sky130_fd_sc_hd__clkbuf_2 _28130_ (.A(_07334_),
    .X(_07335_));
 sky130_fd_sc_hd__a211o_1 _28131_ (.A1(\irq_mask[0] ),
    .A2(_07331_),
    .B1(_07333_),
    .C1(_07335_),
    .X(_01033_));
 sky130_fd_sc_hd__nor2_1 _28132_ (.A(_08744_),
    .B(_07332_),
    .Y(_07336_));
 sky130_fd_sc_hd__clkbuf_2 _28133_ (.A(_07334_),
    .X(_07337_));
 sky130_fd_sc_hd__a211o_1 _28134_ (.A1(_08281_),
    .A2(_07331_),
    .B1(_07336_),
    .C1(_07337_),
    .X(_01034_));
 sky130_fd_sc_hd__nor2_1 _28135_ (.A(_08798_),
    .B(_07332_),
    .Y(_07338_));
 sky130_fd_sc_hd__a211o_1 _28136_ (.A1(\irq_mask[2] ),
    .A2(_07331_),
    .B1(_07338_),
    .C1(_07337_),
    .X(_01035_));
 sky130_fd_sc_hd__nor2_1 _28137_ (.A(_08865_),
    .B(_07332_),
    .Y(_07339_));
 sky130_fd_sc_hd__a211o_1 _28138_ (.A1(\irq_mask[3] ),
    .A2(_07331_),
    .B1(_07339_),
    .C1(_07337_),
    .X(_01036_));
 sky130_fd_sc_hd__clkbuf_2 _28139_ (.A(_07329_),
    .X(_07340_));
 sky130_fd_sc_hd__clkbuf_2 _28140_ (.A(_07340_),
    .X(_07341_));
 sky130_fd_sc_hd__nor2_1 _28141_ (.A(_08934_),
    .B(_07341_),
    .Y(_07342_));
 sky130_fd_sc_hd__a211o_1 _28142_ (.A1(\irq_mask[4] ),
    .A2(_07331_),
    .B1(_07342_),
    .C1(_07337_),
    .X(_01037_));
 sky130_fd_sc_hd__nor2_1 _28143_ (.A(_08978_),
    .B(_07341_),
    .Y(_07343_));
 sky130_fd_sc_hd__a211o_1 _28144_ (.A1(\irq_mask[5] ),
    .A2(_07331_),
    .B1(_07343_),
    .C1(_07337_),
    .X(_01038_));
 sky130_fd_sc_hd__clkbuf_2 _28145_ (.A(_07330_),
    .X(_07344_));
 sky130_fd_sc_hd__nor2_1 _28146_ (.A(_09033_),
    .B(_07341_),
    .Y(_07345_));
 sky130_fd_sc_hd__a211o_1 _28147_ (.A1(\irq_mask[6] ),
    .A2(_07344_),
    .B1(_07345_),
    .C1(_07337_),
    .X(_01039_));
 sky130_fd_sc_hd__nor2_1 _28148_ (.A(_09093_),
    .B(_07341_),
    .Y(_07346_));
 sky130_fd_sc_hd__clkbuf_2 _28149_ (.A(_07334_),
    .X(_07347_));
 sky130_fd_sc_hd__a211o_1 _28150_ (.A1(\irq_mask[7] ),
    .A2(_07344_),
    .B1(_07346_),
    .C1(_07347_),
    .X(_01040_));
 sky130_fd_sc_hd__nor2_1 _28151_ (.A(_09151_),
    .B(_07341_),
    .Y(_07348_));
 sky130_fd_sc_hd__a211o_1 _28152_ (.A1(\irq_mask[8] ),
    .A2(_07344_),
    .B1(_07348_),
    .C1(_07347_),
    .X(_01041_));
 sky130_fd_sc_hd__nor2_1 _28153_ (.A(_09205_),
    .B(_07341_),
    .Y(_07349_));
 sky130_fd_sc_hd__a211o_1 _28154_ (.A1(\irq_mask[9] ),
    .A2(_07344_),
    .B1(_07349_),
    .C1(_07347_),
    .X(_01042_));
 sky130_fd_sc_hd__clkbuf_2 _28155_ (.A(_07340_),
    .X(_07350_));
 sky130_fd_sc_hd__nor2_1 _28156_ (.A(_09245_),
    .B(_07350_),
    .Y(_07351_));
 sky130_fd_sc_hd__a211o_1 _28157_ (.A1(\irq_mask[10] ),
    .A2(_07344_),
    .B1(_07351_),
    .C1(_07347_),
    .X(_01043_));
 sky130_fd_sc_hd__nor2_1 _28158_ (.A(_09282_),
    .B(_07350_),
    .Y(_07352_));
 sky130_fd_sc_hd__a211o_1 _28159_ (.A1(\irq_mask[11] ),
    .A2(_07344_),
    .B1(_07352_),
    .C1(_07347_),
    .X(_01044_));
 sky130_fd_sc_hd__clkbuf_2 _28160_ (.A(_07340_),
    .X(_07353_));
 sky130_fd_sc_hd__nor2_1 _28161_ (.A(_09332_),
    .B(_07350_),
    .Y(_07354_));
 sky130_fd_sc_hd__a211o_1 _28162_ (.A1(\irq_mask[12] ),
    .A2(_07353_),
    .B1(_07354_),
    .C1(_07347_),
    .X(_01045_));
 sky130_fd_sc_hd__nor2_1 _28163_ (.A(_09372_),
    .B(_07350_),
    .Y(_07355_));
 sky130_fd_sc_hd__clkbuf_2 _28164_ (.A(_07334_),
    .X(_07356_));
 sky130_fd_sc_hd__a211o_1 _28165_ (.A1(\irq_mask[13] ),
    .A2(_07353_),
    .B1(_07355_),
    .C1(_07356_),
    .X(_01046_));
 sky130_fd_sc_hd__nor2_1 _28166_ (.A(_09414_),
    .B(_07350_),
    .Y(_07357_));
 sky130_fd_sc_hd__a211o_1 _28167_ (.A1(\irq_mask[14] ),
    .A2(_07353_),
    .B1(_07357_),
    .C1(_07356_),
    .X(_01047_));
 sky130_fd_sc_hd__nor2_1 _28168_ (.A(_09453_),
    .B(_07350_),
    .Y(_07358_));
 sky130_fd_sc_hd__a211o_1 _28169_ (.A1(\irq_mask[15] ),
    .A2(_07353_),
    .B1(_07358_),
    .C1(_07356_),
    .X(_01048_));
 sky130_fd_sc_hd__clkbuf_2 _28170_ (.A(_07340_),
    .X(_07359_));
 sky130_fd_sc_hd__nor2_1 _28171_ (.A(_09507_),
    .B(_07359_),
    .Y(_07360_));
 sky130_fd_sc_hd__a211o_1 _28172_ (.A1(\irq_mask[16] ),
    .A2(_07353_),
    .B1(_07360_),
    .C1(_07356_),
    .X(_01049_));
 sky130_fd_sc_hd__nor2_1 _28173_ (.A(_09545_),
    .B(_07359_),
    .Y(_07361_));
 sky130_fd_sc_hd__a211o_1 _28174_ (.A1(\irq_mask[17] ),
    .A2(_07353_),
    .B1(_07361_),
    .C1(_07356_),
    .X(_01050_));
 sky130_fd_sc_hd__clkbuf_2 _28175_ (.A(_07340_),
    .X(_07362_));
 sky130_fd_sc_hd__nor2_1 _28176_ (.A(_09589_),
    .B(_07359_),
    .Y(_07363_));
 sky130_fd_sc_hd__a211o_1 _28177_ (.A1(\irq_mask[18] ),
    .A2(_07362_),
    .B1(_07363_),
    .C1(_07356_),
    .X(_01051_));
 sky130_fd_sc_hd__nor2_1 _28178_ (.A(_09626_),
    .B(_07359_),
    .Y(_07364_));
 sky130_fd_sc_hd__clkbuf_2 _28179_ (.A(_07334_),
    .X(_07365_));
 sky130_fd_sc_hd__a211o_1 _28180_ (.A1(\irq_mask[19] ),
    .A2(_07362_),
    .B1(_07364_),
    .C1(_07365_),
    .X(_01052_));
 sky130_fd_sc_hd__nor2_1 _28181_ (.A(_09667_),
    .B(_07359_),
    .Y(_07366_));
 sky130_fd_sc_hd__a211o_1 _28182_ (.A1(\irq_mask[20] ),
    .A2(_07362_),
    .B1(_07366_),
    .C1(_07365_),
    .X(_01053_));
 sky130_fd_sc_hd__nor2_1 _28183_ (.A(_09704_),
    .B(_07359_),
    .Y(_07367_));
 sky130_fd_sc_hd__a211o_1 _28184_ (.A1(\irq_mask[21] ),
    .A2(_07362_),
    .B1(_07367_),
    .C1(_07365_),
    .X(_01054_));
 sky130_fd_sc_hd__clkbuf_2 _28185_ (.A(_07329_),
    .X(_07368_));
 sky130_fd_sc_hd__nor2_1 _28186_ (.A(_09744_),
    .B(_07368_),
    .Y(_07369_));
 sky130_fd_sc_hd__a211o_1 _28187_ (.A1(\irq_mask[22] ),
    .A2(_07362_),
    .B1(_07369_),
    .C1(_07365_),
    .X(_01055_));
 sky130_fd_sc_hd__nor2_1 _28188_ (.A(_09781_),
    .B(_07368_),
    .Y(_07370_));
 sky130_fd_sc_hd__a211o_1 _28189_ (.A1(\irq_mask[23] ),
    .A2(_07362_),
    .B1(_07370_),
    .C1(_07365_),
    .X(_01056_));
 sky130_fd_sc_hd__clkbuf_2 _28190_ (.A(_07340_),
    .X(_07371_));
 sky130_fd_sc_hd__nor2_1 _28191_ (.A(_09821_),
    .B(_07368_),
    .Y(_07372_));
 sky130_fd_sc_hd__a211o_1 _28192_ (.A1(\irq_mask[24] ),
    .A2(_07371_),
    .B1(_07372_),
    .C1(_07365_),
    .X(_01057_));
 sky130_fd_sc_hd__nor2_1 _28193_ (.A(_09855_),
    .B(_07368_),
    .Y(_07373_));
 sky130_fd_sc_hd__clkbuf_2 _28194_ (.A(_06200_),
    .X(_07374_));
 sky130_fd_sc_hd__a211o_1 _28195_ (.A1(\irq_mask[25] ),
    .A2(_07371_),
    .B1(_07373_),
    .C1(_07374_),
    .X(_01058_));
 sky130_fd_sc_hd__nor2_1 _28196_ (.A(_09888_),
    .B(_07368_),
    .Y(_07375_));
 sky130_fd_sc_hd__a211o_1 _28197_ (.A1(\irq_mask[26] ),
    .A2(_07371_),
    .B1(_07375_),
    .C1(_07374_),
    .X(_01059_));
 sky130_fd_sc_hd__nor2_1 _28198_ (.A(_09929_),
    .B(_07368_),
    .Y(_07376_));
 sky130_fd_sc_hd__a211o_1 _28199_ (.A1(\irq_mask[27] ),
    .A2(_07371_),
    .B1(_07376_),
    .C1(_07374_),
    .X(_01060_));
 sky130_fd_sc_hd__nor2_1 _28200_ (.A(_09966_),
    .B(_07330_),
    .Y(_07377_));
 sky130_fd_sc_hd__a211o_1 _28201_ (.A1(\irq_mask[28] ),
    .A2(_07371_),
    .B1(_07377_),
    .C1(_07374_),
    .X(_01061_));
 sky130_fd_sc_hd__nor2_1 _28202_ (.A(_10003_),
    .B(_07330_),
    .Y(_07378_));
 sky130_fd_sc_hd__a211o_1 _28203_ (.A1(\irq_mask[29] ),
    .A2(_07371_),
    .B1(_07378_),
    .C1(_07374_),
    .X(_01062_));
 sky130_fd_sc_hd__nor2_1 _28204_ (.A(_10040_),
    .B(_07330_),
    .Y(_07379_));
 sky130_fd_sc_hd__a211o_1 _28205_ (.A1(\irq_mask[30] ),
    .A2(_07332_),
    .B1(_07379_),
    .C1(_07374_),
    .X(_01063_));
 sky130_fd_sc_hd__nor2_1 _28206_ (.A(_10077_),
    .B(_07330_),
    .Y(_07380_));
 sky130_fd_sc_hd__a211o_1 _28207_ (.A1(\irq_mask[31] ),
    .A2(_07332_),
    .B1(_07380_),
    .C1(_06201_),
    .X(_01064_));
 sky130_fd_sc_hd__and2_2 _28208_ (.A(_08328_),
    .B(_08538_),
    .X(_07381_));
 sky130_fd_sc_hd__clkbuf_2 _28209_ (.A(_07381_),
    .X(_07382_));
 sky130_fd_sc_hd__nand2_1 _28210_ (.A(_08146_),
    .B(_08538_),
    .Y(_07383_));
 sky130_fd_sc_hd__clkbuf_2 _28211_ (.A(_07383_),
    .X(_07384_));
 sky130_fd_sc_hd__buf_2 _28212_ (.A(is_slli_srli_srai),
    .X(_07385_));
 sky130_fd_sc_hd__mux2_1 _28213_ (.A0(_08668_),
    .A1(_08554_),
    .S(_07385_),
    .X(_07386_));
 sky130_fd_sc_hd__nor2_1 _28214_ (.A(_08902_),
    .B(_07386_),
    .Y(_07387_));
 sky130_fd_sc_hd__a211o_1 _28215_ (.A1(_08518_),
    .A2(_08635_),
    .B1(_07384_),
    .C1(_07387_),
    .X(_07388_));
 sky130_fd_sc_hd__o21ai_1 _28216_ (.A1(_08470_),
    .A2(_07382_),
    .B1(_07388_),
    .Y(_01065_));
 sky130_fd_sc_hd__buf_2 _28217_ (.A(_07384_),
    .X(_07389_));
 sky130_fd_sc_hd__mux2_1 _28218_ (.A0(_08762_),
    .A1(_08546_),
    .S(_07385_),
    .X(_07390_));
 sky130_fd_sc_hd__or2_1 _28219_ (.A(_09520_),
    .B(_07390_),
    .X(_07391_));
 sky130_fd_sc_hd__a21oi_1 _28220_ (.A1(_08518_),
    .A2(_08744_),
    .B1(_07389_),
    .Y(_07392_));
 sky130_fd_sc_hd__a22o_1 _28221_ (.A1(_10108_),
    .A2(_07389_),
    .B1(_07391_),
    .B2(_07392_),
    .X(_01066_));
 sky130_fd_sc_hd__mux2_1 _28222_ (.A0(\decoded_imm[2] ),
    .A1(\decoded_imm_uj[2] ),
    .S(_07385_),
    .X(_07393_));
 sky130_fd_sc_hd__or2_1 _28223_ (.A(_09600_),
    .B(_07393_),
    .X(_07394_));
 sky130_fd_sc_hd__clkbuf_2 _28224_ (.A(_07383_),
    .X(_07395_));
 sky130_fd_sc_hd__a21oi_1 _28225_ (.A1(_08518_),
    .A2(_08798_),
    .B1(_07395_),
    .Y(_07396_));
 sky130_fd_sc_hd__a22o_1 _28226_ (.A1(_10273_),
    .A2(_07389_),
    .B1(_07394_),
    .B2(_07396_),
    .X(_01067_));
 sky130_fd_sc_hd__buf_2 _28227_ (.A(_04768_),
    .X(_07397_));
 sky130_fd_sc_hd__mux2_1 _28228_ (.A0(\decoded_imm[3] ),
    .A1(\decoded_imm_uj[3] ),
    .S(_07385_),
    .X(_07398_));
 sky130_fd_sc_hd__or2_1 _28229_ (.A(_09600_),
    .B(_07398_),
    .X(_07399_));
 sky130_fd_sc_hd__a21oi_1 _28230_ (.A1(_08518_),
    .A2(_08865_),
    .B1(_07395_),
    .Y(_07400_));
 sky130_fd_sc_hd__a22o_1 _28231_ (.A1(_07397_),
    .A2(_07389_),
    .B1(_07399_),
    .B2(_07400_),
    .X(_01068_));
 sky130_fd_sc_hd__mux2_1 _28232_ (.A0(\decoded_imm[4] ),
    .A1(\decoded_imm_uj[4] ),
    .S(_07385_),
    .X(_07401_));
 sky130_fd_sc_hd__or2_1 _28233_ (.A(_09600_),
    .B(_07401_),
    .X(_07402_));
 sky130_fd_sc_hd__a21oi_1 _28234_ (.A1(_08518_),
    .A2(_08934_),
    .B1(_07395_),
    .Y(_07403_));
 sky130_fd_sc_hd__a22o_1 _28235_ (.A1(_04756_),
    .A2(_07389_),
    .B1(_07402_),
    .B2(_07403_),
    .X(_01069_));
 sky130_fd_sc_hd__clkbuf_2 _28236_ (.A(_07382_),
    .X(_07404_));
 sky130_vsdinv _28237_ (.A(_08978_),
    .Y(_07405_));
 sky130_fd_sc_hd__nor2_1 _28238_ (.A(_08287_),
    .B(is_slli_srli_srai),
    .Y(_07406_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28239_ (.A(_07406_),
    .X(_07407_));
 sky130_fd_sc_hd__clkbuf_2 _28240_ (.A(_07407_),
    .X(_07408_));
 sky130_fd_sc_hd__a221o_1 _28241_ (.A1(_09291_),
    .A2(_07405_),
    .B1(_07408_),
    .B2(\decoded_imm[5] ),
    .C1(_07395_),
    .X(_07409_));
 sky130_fd_sc_hd__o21a_1 _28242_ (.A1(_10277_),
    .A2(_07404_),
    .B1(_07409_),
    .X(_01070_));
 sky130_vsdinv _28243_ (.A(_09033_),
    .Y(_07410_));
 sky130_fd_sc_hd__a221o_1 _28244_ (.A1(_09291_),
    .A2(_07410_),
    .B1(_07408_),
    .B2(\decoded_imm[6] ),
    .C1(_07395_),
    .X(_07411_));
 sky130_fd_sc_hd__o21a_1 _28245_ (.A1(_10279_),
    .A2(_07404_),
    .B1(_07411_),
    .X(_01071_));
 sky130_vsdinv _28246_ (.A(_09093_),
    .Y(_07412_));
 sky130_fd_sc_hd__a221o_1 _28247_ (.A1(_09291_),
    .A2(_07412_),
    .B1(_07408_),
    .B2(\decoded_imm[7] ),
    .C1(_07395_),
    .X(_07413_));
 sky130_fd_sc_hd__o21a_1 _28248_ (.A1(_10280_),
    .A2(_07404_),
    .B1(_07413_),
    .X(_01072_));
 sky130_vsdinv _28249_ (.A(_09151_),
    .Y(_07414_));
 sky130_fd_sc_hd__clkbuf_2 _28250_ (.A(_07384_),
    .X(_07415_));
 sky130_fd_sc_hd__a221o_1 _28251_ (.A1(_09291_),
    .A2(_07414_),
    .B1(_07408_),
    .B2(\decoded_imm[8] ),
    .C1(_07415_),
    .X(_07416_));
 sky130_fd_sc_hd__o21a_1 _28252_ (.A1(_08484_),
    .A2(_07404_),
    .B1(_07416_),
    .X(_01073_));
 sky130_vsdinv _28253_ (.A(_09205_),
    .Y(_07417_));
 sky130_fd_sc_hd__a221o_1 _28254_ (.A1(_09291_),
    .A2(_07417_),
    .B1(_07408_),
    .B2(\decoded_imm[9] ),
    .C1(_07415_),
    .X(_07418_));
 sky130_fd_sc_hd__o21a_1 _28255_ (.A1(_10158_),
    .A2(_07404_),
    .B1(_07418_),
    .X(_01074_));
 sky130_fd_sc_hd__clkbuf_2 _28256_ (.A(_08517_),
    .X(_07419_));
 sky130_vsdinv _28257_ (.A(_09245_),
    .Y(_07420_));
 sky130_fd_sc_hd__a221o_1 _28258_ (.A1(_07419_),
    .A2(_07420_),
    .B1(_07408_),
    .B2(_09219_),
    .C1(_07415_),
    .X(_07421_));
 sky130_fd_sc_hd__o21a_1 _28259_ (.A1(_10164_),
    .A2(_07404_),
    .B1(_07421_),
    .X(_01075_));
 sky130_fd_sc_hd__clkbuf_2 _28260_ (.A(_07382_),
    .X(_07422_));
 sky130_vsdinv _28261_ (.A(_09282_),
    .Y(_07423_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28262_ (.A(_07407_),
    .X(_07424_));
 sky130_fd_sc_hd__a221o_1 _28263_ (.A1(_07419_),
    .A2(_07423_),
    .B1(_07424_),
    .B2(\decoded_imm[11] ),
    .C1(_07415_),
    .X(_07425_));
 sky130_fd_sc_hd__o21a_1 _28264_ (.A1(_08413_),
    .A2(_07422_),
    .B1(_07425_),
    .X(_01076_));
 sky130_vsdinv _28265_ (.A(_09332_),
    .Y(_07426_));
 sky130_fd_sc_hd__a221o_1 _28266_ (.A1(_07419_),
    .A2(_07426_),
    .B1(_07424_),
    .B2(_09305_),
    .C1(_07415_),
    .X(_07427_));
 sky130_fd_sc_hd__o21a_1 _28267_ (.A1(_08343_),
    .A2(_07422_),
    .B1(_07427_),
    .X(_01077_));
 sky130_vsdinv _28268_ (.A(_09372_),
    .Y(_07428_));
 sky130_fd_sc_hd__a221o_1 _28269_ (.A1(_07419_),
    .A2(_07428_),
    .B1(_07424_),
    .B2(\decoded_imm[13] ),
    .C1(_07415_),
    .X(_07429_));
 sky130_fd_sc_hd__o21a_1 _28270_ (.A1(_08347_),
    .A2(_07422_),
    .B1(_07429_),
    .X(_01078_));
 sky130_vsdinv _28271_ (.A(_09414_),
    .Y(_07430_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28272_ (.A(_07384_),
    .X(_07431_));
 sky130_fd_sc_hd__a221o_1 _28273_ (.A1(_07419_),
    .A2(_07430_),
    .B1(_07424_),
    .B2(\decoded_imm[14] ),
    .C1(_07431_),
    .X(_07432_));
 sky130_fd_sc_hd__o21a_1 _28274_ (.A1(_08419_),
    .A2(_07422_),
    .B1(_07432_),
    .X(_01079_));
 sky130_vsdinv _28275_ (.A(_09453_),
    .Y(_07433_));
 sky130_fd_sc_hd__a221o_1 _28276_ (.A1(_07419_),
    .A2(_07433_),
    .B1(_07424_),
    .B2(\decoded_imm[15] ),
    .C1(_07431_),
    .X(_07434_));
 sky130_fd_sc_hd__o21a_1 _28277_ (.A1(_10188_),
    .A2(_07422_),
    .B1(_07434_),
    .X(_01080_));
 sky130_fd_sc_hd__clkbuf_2 _28278_ (.A(_08771_),
    .X(_07435_));
 sky130_vsdinv _28279_ (.A(_09507_),
    .Y(_07436_));
 sky130_fd_sc_hd__a221o_1 _28280_ (.A1(_07435_),
    .A2(_07436_),
    .B1(_07424_),
    .B2(\decoded_imm[16] ),
    .C1(_07431_),
    .X(_07437_));
 sky130_fd_sc_hd__o21a_1 _28281_ (.A1(net306),
    .A2(_07422_),
    .B1(_07437_),
    .X(_01081_));
 sky130_fd_sc_hd__clkbuf_2 _28282_ (.A(_07381_),
    .X(_07438_));
 sky130_vsdinv _28283_ (.A(_09545_),
    .Y(_07439_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28284_ (.A(_07407_),
    .X(_07440_));
 sky130_fd_sc_hd__a221o_1 _28285_ (.A1(_07435_),
    .A2(_07439_),
    .B1(_07440_),
    .B2(\decoded_imm[17] ),
    .C1(_07431_),
    .X(_07441_));
 sky130_fd_sc_hd__o21a_1 _28286_ (.A1(_08383_),
    .A2(_07438_),
    .B1(_07441_),
    .X(_01082_));
 sky130_vsdinv _28287_ (.A(_09589_),
    .Y(_07442_));
 sky130_fd_sc_hd__a221o_1 _28288_ (.A1(_07435_),
    .A2(_07442_),
    .B1(_07440_),
    .B2(\decoded_imm[18] ),
    .C1(_07431_),
    .X(_07443_));
 sky130_fd_sc_hd__o21a_1 _28289_ (.A1(net308),
    .A2(_07438_),
    .B1(_07443_),
    .X(_01083_));
 sky130_vsdinv _28290_ (.A(_09626_),
    .Y(_07444_));
 sky130_fd_sc_hd__a221o_1 _28291_ (.A1(_07435_),
    .A2(_07444_),
    .B1(_07440_),
    .B2(\decoded_imm[19] ),
    .C1(_07431_),
    .X(_07445_));
 sky130_fd_sc_hd__o21a_1 _28292_ (.A1(_08375_),
    .A2(_07438_),
    .B1(_07445_),
    .X(_01084_));
 sky130_vsdinv _28293_ (.A(_09667_),
    .Y(_07446_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28294_ (.A(_07384_),
    .X(_07447_));
 sky130_fd_sc_hd__a221o_1 _28295_ (.A1(_07435_),
    .A2(_07446_),
    .B1(_07440_),
    .B2(\decoded_imm[20] ),
    .C1(_07447_),
    .X(_07448_));
 sky130_fd_sc_hd__o21a_1 _28296_ (.A1(net311),
    .A2(_07438_),
    .B1(_07448_),
    .X(_01085_));
 sky130_vsdinv _28297_ (.A(_09704_),
    .Y(_07449_));
 sky130_fd_sc_hd__a221o_1 _28298_ (.A1(_07435_),
    .A2(_07449_),
    .B1(_07440_),
    .B2(\decoded_imm[21] ),
    .C1(_07447_),
    .X(_07450_));
 sky130_fd_sc_hd__o21a_1 _28299_ (.A1(_08364_),
    .A2(_07438_),
    .B1(_07450_),
    .X(_01086_));
 sky130_fd_sc_hd__clkbuf_2 _28300_ (.A(_08771_),
    .X(_07451_));
 sky130_vsdinv _28301_ (.A(_09744_),
    .Y(_07452_));
 sky130_fd_sc_hd__a221o_1 _28302_ (.A1(_07451_),
    .A2(_07452_),
    .B1(_07440_),
    .B2(\decoded_imm[22] ),
    .C1(_07447_),
    .X(_07453_));
 sky130_fd_sc_hd__o21a_1 _28303_ (.A1(net313),
    .A2(_07438_),
    .B1(_07453_),
    .X(_01087_));
 sky130_fd_sc_hd__clkbuf_2 _28304_ (.A(_07381_),
    .X(_07454_));
 sky130_vsdinv _28305_ (.A(_09781_),
    .Y(_07455_));
 sky130_fd_sc_hd__clkbuf_2 _28306_ (.A(_07406_),
    .X(_07456_));
 sky130_fd_sc_hd__a221o_1 _28307_ (.A1(_07451_),
    .A2(_07455_),
    .B1(_07456_),
    .B2(_09751_),
    .C1(_07447_),
    .X(_07457_));
 sky130_fd_sc_hd__o21a_1 _28308_ (.A1(_08369_),
    .A2(_07454_),
    .B1(_07457_),
    .X(_01088_));
 sky130_vsdinv _28309_ (.A(_09821_),
    .Y(_07458_));
 sky130_fd_sc_hd__a221o_1 _28310_ (.A1(_07451_),
    .A2(_07458_),
    .B1(_07456_),
    .B2(\decoded_imm[24] ),
    .C1(_07447_),
    .X(_07459_));
 sky130_fd_sc_hd__o21a_1 _28311_ (.A1(net315),
    .A2(_07454_),
    .B1(_07459_),
    .X(_01089_));
 sky130_vsdinv _28312_ (.A(_09855_),
    .Y(_07460_));
 sky130_fd_sc_hd__a221o_1 _28313_ (.A1(_07451_),
    .A2(_07460_),
    .B1(_07456_),
    .B2(\decoded_imm[25] ),
    .C1(_07447_),
    .X(_07461_));
 sky130_fd_sc_hd__o21a_1 _28314_ (.A1(_08427_),
    .A2(_07454_),
    .B1(_07461_),
    .X(_01090_));
 sky130_vsdinv _28315_ (.A(_09888_),
    .Y(_07462_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28316_ (.A(_07384_),
    .X(_07463_));
 sky130_fd_sc_hd__a221o_1 _28317_ (.A1(_07451_),
    .A2(_07462_),
    .B1(_07456_),
    .B2(\decoded_imm[26] ),
    .C1(_07463_),
    .X(_07464_));
 sky130_fd_sc_hd__o21a_1 _28318_ (.A1(net317),
    .A2(_07454_),
    .B1(_07464_),
    .X(_01091_));
 sky130_vsdinv _28319_ (.A(_09929_),
    .Y(_07465_));
 sky130_fd_sc_hd__a221o_1 _28320_ (.A1(_07451_),
    .A2(_07465_),
    .B1(_07456_),
    .B2(\decoded_imm[27] ),
    .C1(_07463_),
    .X(_07466_));
 sky130_fd_sc_hd__o21a_1 _28321_ (.A1(_08436_),
    .A2(_07454_),
    .B1(_07466_),
    .X(_01092_));
 sky130_vsdinv _28322_ (.A(_09966_),
    .Y(_07467_));
 sky130_fd_sc_hd__a221o_1 _28323_ (.A1(_09520_),
    .A2(_07467_),
    .B1(_07456_),
    .B2(\decoded_imm[28] ),
    .C1(_07463_),
    .X(_07468_));
 sky130_fd_sc_hd__o21a_1 _28324_ (.A1(_08479_),
    .A2(_07454_),
    .B1(_07468_),
    .X(_01093_));
 sky130_vsdinv _28325_ (.A(_10003_),
    .Y(_07469_));
 sky130_fd_sc_hd__a221o_1 _28326_ (.A1(_09520_),
    .A2(_07469_),
    .B1(_07407_),
    .B2(\decoded_imm[29] ),
    .C1(_07463_),
    .X(_07470_));
 sky130_fd_sc_hd__o21a_1 _28327_ (.A1(_08398_),
    .A2(_07382_),
    .B1(_07470_),
    .X(_01094_));
 sky130_vsdinv _28328_ (.A(_10040_),
    .Y(_07471_));
 sky130_fd_sc_hd__a221o_1 _28329_ (.A1(_09520_),
    .A2(_07471_),
    .B1(_07407_),
    .B2(\decoded_imm[30] ),
    .C1(_07463_),
    .X(_07472_));
 sky130_fd_sc_hd__o21a_1 _28330_ (.A1(_08487_),
    .A2(_07382_),
    .B1(_07472_),
    .X(_01095_));
 sky130_vsdinv _28331_ (.A(_10077_),
    .Y(_07473_));
 sky130_fd_sc_hd__a221o_1 _28332_ (.A1(_09520_),
    .A2(_07473_),
    .B1(_07407_),
    .B2(\decoded_imm[31] ),
    .C1(_07463_),
    .X(_07474_));
 sky130_fd_sc_hd__o21a_1 _28333_ (.A1(_10260_),
    .A2(_07382_),
    .B1(_07474_),
    .X(_01096_));
 sky130_fd_sc_hd__clkbuf_2 _28334_ (.A(_10306_),
    .X(_07475_));
 sky130_fd_sc_hd__clkbuf_2 _28335_ (.A(_07475_),
    .X(_07476_));
 sky130_fd_sc_hd__clkbuf_2 _28336_ (.A(_10307_),
    .X(_07477_));
 sky130_fd_sc_hd__clkbuf_2 _28337_ (.A(_07477_),
    .X(_07478_));
 sky130_fd_sc_hd__or4_2 _28338_ (.A(\timer[29] ),
    .B(\timer[28] ),
    .C(\timer[31] ),
    .D(\timer[30] ),
    .X(_07479_));
 sky130_fd_sc_hd__or4_2 _28339_ (.A(\timer[21] ),
    .B(\timer[20] ),
    .C(\timer[23] ),
    .D(\timer[22] ),
    .X(_07480_));
 sky130_fd_sc_hd__or4_2 _28340_ (.A(\timer[5] ),
    .B(\timer[4] ),
    .C(\timer[7] ),
    .D(\timer[6] ),
    .X(_07481_));
 sky130_fd_sc_hd__or4_1 _28341_ (.A(\timer[13] ),
    .B(\timer[12] ),
    .C(\timer[15] ),
    .D(\timer[14] ),
    .X(_07482_));
 sky130_fd_sc_hd__or4_1 _28342_ (.A(\timer[3] ),
    .B(\timer[2] ),
    .C(\timer[11] ),
    .D(_09247_),
    .X(_07483_));
 sky130_fd_sc_hd__or4_1 _28343_ (.A(\timer[19] ),
    .B(\timer[18] ),
    .C(\timer[27] ),
    .D(\timer[26] ),
    .X(_07484_));
 sky130_fd_sc_hd__or4b_1 _28344_ (.A(\timer[1] ),
    .B(\timer[9] ),
    .C(\timer[8] ),
    .D_N(\timer[0] ),
    .X(_07485_));
 sky130_fd_sc_hd__or4_1 _28345_ (.A(\timer[17] ),
    .B(\timer[16] ),
    .C(\timer[25] ),
    .D(\timer[24] ),
    .X(_07486_));
 sky130_fd_sc_hd__or4_1 _28346_ (.A(_07483_),
    .B(_07484_),
    .C(_07485_),
    .D(_07486_),
    .X(_07487_));
 sky130_fd_sc_hd__or4_1 _28347_ (.A(_07480_),
    .B(_07481_),
    .C(_07482_),
    .D(_07487_),
    .X(_07488_));
 sky130_fd_sc_hd__nor2_1 _28348_ (.A(_07479_),
    .B(_07488_),
    .Y(_07489_));
 sky130_fd_sc_hd__or3_1 _28349_ (.A(\irq_pending[0] ),
    .B(net1),
    .C(_07489_),
    .X(_07490_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28350_ (.A(_07327_),
    .X(_07491_));
 sky130_fd_sc_hd__o311a_1 _28351_ (.A1(_07476_),
    .A2(\irq_mask[0] ),
    .A3(_07478_),
    .B1(_07490_),
    .C1(_07491_),
    .X(_01097_));
 sky130_fd_sc_hd__o32a_1 _28352_ (.A1(_07475_),
    .A2(_08281_),
    .A3(_07477_),
    .B1(net12),
    .B2(\irq_pending[1] ),
    .X(_07492_));
 sky130_fd_sc_hd__nor4_1 _28353_ (.A(_08281_),
    .B(_08186_),
    .C(_08282_),
    .D(_08319_),
    .Y(_07493_));
 sky130_fd_sc_hd__o21a_1 _28354_ (.A1(_07492_),
    .A2(_07493_),
    .B1(_06130_),
    .X(_01098_));
 sky130_fd_sc_hd__or2_1 _28355_ (.A(\irq_pending[3] ),
    .B(net26),
    .X(_07494_));
 sky130_fd_sc_hd__o311a_1 _28356_ (.A1(_07476_),
    .A2(\irq_mask[3] ),
    .A3(_07478_),
    .B1(_07494_),
    .C1(_07491_),
    .X(_01099_));
 sky130_fd_sc_hd__or2_1 _28357_ (.A(\irq_pending[4] ),
    .B(net27),
    .X(_07495_));
 sky130_fd_sc_hd__o311a_1 _28358_ (.A1(_07476_),
    .A2(\irq_mask[4] ),
    .A3(_07478_),
    .B1(_07495_),
    .C1(_07491_),
    .X(_01100_));
 sky130_fd_sc_hd__or2_1 _28359_ (.A(\irq_pending[5] ),
    .B(net28),
    .X(_07496_));
 sky130_fd_sc_hd__o311a_1 _28360_ (.A1(_07476_),
    .A2(\irq_mask[5] ),
    .A3(_07478_),
    .B1(_07496_),
    .C1(_07491_),
    .X(_01101_));
 sky130_fd_sc_hd__or2_1 _28361_ (.A(\irq_pending[6] ),
    .B(net29),
    .X(_07497_));
 sky130_fd_sc_hd__o311a_1 _28362_ (.A1(_07476_),
    .A2(\irq_mask[6] ),
    .A3(_07478_),
    .B1(_07497_),
    .C1(_07491_),
    .X(_01102_));
 sky130_fd_sc_hd__or2_1 _28363_ (.A(\irq_pending[7] ),
    .B(net30),
    .X(_07498_));
 sky130_fd_sc_hd__o311a_1 _28364_ (.A1(_07476_),
    .A2(\irq_mask[7] ),
    .A3(_07478_),
    .B1(_07498_),
    .C1(_07491_),
    .X(_01103_));
 sky130_fd_sc_hd__clkbuf_2 _28365_ (.A(_07475_),
    .X(_07499_));
 sky130_fd_sc_hd__clkbuf_2 _28366_ (.A(_07477_),
    .X(_07500_));
 sky130_fd_sc_hd__or2_1 _28367_ (.A(\irq_pending[8] ),
    .B(net31),
    .X(_07501_));
 sky130_fd_sc_hd__clkbuf_2 _28368_ (.A(_07327_),
    .X(_07502_));
 sky130_fd_sc_hd__o311a_1 _28369_ (.A1(_07499_),
    .A2(net449),
    .A3(_07500_),
    .B1(_07501_),
    .C1(_07502_),
    .X(_01104_));
 sky130_fd_sc_hd__or2_1 _28370_ (.A(\irq_pending[9] ),
    .B(net32),
    .X(_07503_));
 sky130_fd_sc_hd__o311a_1 _28371_ (.A1(_07499_),
    .A2(net440),
    .A3(_07500_),
    .B1(_07503_),
    .C1(_07502_),
    .X(_01105_));
 sky130_fd_sc_hd__or2_1 _28372_ (.A(\irq_pending[10] ),
    .B(net2),
    .X(_07504_));
 sky130_fd_sc_hd__o311a_1 _28373_ (.A1(_07499_),
    .A2(net448),
    .A3(_07500_),
    .B1(_07504_),
    .C1(_07502_),
    .X(_01106_));
 sky130_fd_sc_hd__or2_1 _28374_ (.A(\irq_pending[11] ),
    .B(net3),
    .X(_07505_));
 sky130_fd_sc_hd__o311a_1 _28375_ (.A1(_07499_),
    .A2(net458),
    .A3(_07500_),
    .B1(_07505_),
    .C1(_07502_),
    .X(_01107_));
 sky130_fd_sc_hd__or2_1 _28376_ (.A(\irq_pending[12] ),
    .B(net4),
    .X(_07506_));
 sky130_fd_sc_hd__o311a_1 _28377_ (.A1(_07499_),
    .A2(net452),
    .A3(_07500_),
    .B1(_07506_),
    .C1(_07502_),
    .X(_01108_));
 sky130_fd_sc_hd__or2_1 _28378_ (.A(\irq_pending[13] ),
    .B(net5),
    .X(_07507_));
 sky130_fd_sc_hd__o311a_1 _28379_ (.A1(_07499_),
    .A2(\irq_mask[13] ),
    .A3(_07500_),
    .B1(_07507_),
    .C1(_07502_),
    .X(_01109_));
 sky130_fd_sc_hd__clkbuf_2 _28380_ (.A(_07475_),
    .X(_07508_));
 sky130_fd_sc_hd__clkbuf_2 _28381_ (.A(_07477_),
    .X(_07509_));
 sky130_fd_sc_hd__or2_1 _28382_ (.A(\irq_pending[14] ),
    .B(net6),
    .X(_07510_));
 sky130_fd_sc_hd__clkbuf_2 _28383_ (.A(_07327_),
    .X(_07511_));
 sky130_fd_sc_hd__o311a_1 _28384_ (.A1(_07508_),
    .A2(\irq_mask[14] ),
    .A3(_07509_),
    .B1(_07510_),
    .C1(_07511_),
    .X(_01110_));
 sky130_fd_sc_hd__or2_1 _28385_ (.A(\irq_pending[15] ),
    .B(net7),
    .X(_07512_));
 sky130_fd_sc_hd__o311a_1 _28386_ (.A1(_07508_),
    .A2(\irq_mask[15] ),
    .A3(_07509_),
    .B1(_07512_),
    .C1(_07511_),
    .X(_01111_));
 sky130_fd_sc_hd__or2_1 _28387_ (.A(\irq_pending[16] ),
    .B(net8),
    .X(_07513_));
 sky130_fd_sc_hd__o311a_1 _28388_ (.A1(_07508_),
    .A2(\irq_mask[16] ),
    .A3(_07509_),
    .B1(_07513_),
    .C1(_07511_),
    .X(_01112_));
 sky130_fd_sc_hd__or2_1 _28389_ (.A(\irq_pending[17] ),
    .B(net9),
    .X(_07514_));
 sky130_fd_sc_hd__o311a_1 _28390_ (.A1(_07508_),
    .A2(\irq_mask[17] ),
    .A3(_07509_),
    .B1(_07514_),
    .C1(_07511_),
    .X(_01113_));
 sky130_fd_sc_hd__or2_1 _28391_ (.A(\irq_pending[18] ),
    .B(net10),
    .X(_07515_));
 sky130_fd_sc_hd__o311a_1 _28392_ (.A1(_07508_),
    .A2(\irq_mask[18] ),
    .A3(_07509_),
    .B1(_07515_),
    .C1(_07511_),
    .X(_01114_));
 sky130_fd_sc_hd__or2_1 _28393_ (.A(\irq_pending[19] ),
    .B(net11),
    .X(_07516_));
 sky130_fd_sc_hd__o311a_1 _28394_ (.A1(_07508_),
    .A2(\irq_mask[19] ),
    .A3(_07509_),
    .B1(_07516_),
    .C1(_07511_),
    .X(_01115_));
 sky130_fd_sc_hd__clkbuf_2 _28395_ (.A(_07475_),
    .X(_07517_));
 sky130_fd_sc_hd__clkbuf_2 _28396_ (.A(_07477_),
    .X(_07518_));
 sky130_fd_sc_hd__or2_1 _28397_ (.A(\irq_pending[20] ),
    .B(net13),
    .X(_07519_));
 sky130_fd_sc_hd__clkbuf_2 _28398_ (.A(_07327_),
    .X(_07520_));
 sky130_fd_sc_hd__o311a_1 _28399_ (.A1(_07517_),
    .A2(\irq_mask[20] ),
    .A3(_07518_),
    .B1(_07519_),
    .C1(_07520_),
    .X(_01116_));
 sky130_fd_sc_hd__or2_1 _28400_ (.A(\irq_pending[21] ),
    .B(net14),
    .X(_07521_));
 sky130_fd_sc_hd__o311a_1 _28401_ (.A1(_07517_),
    .A2(\irq_mask[21] ),
    .A3(_07518_),
    .B1(_07521_),
    .C1(_07520_),
    .X(_01117_));
 sky130_fd_sc_hd__or2_1 _28402_ (.A(\irq_pending[22] ),
    .B(net15),
    .X(_07522_));
 sky130_fd_sc_hd__o311a_1 _28403_ (.A1(_07517_),
    .A2(\irq_mask[22] ),
    .A3(_07518_),
    .B1(_07522_),
    .C1(_07520_),
    .X(_01118_));
 sky130_fd_sc_hd__or2_1 _28404_ (.A(\irq_pending[23] ),
    .B(net16),
    .X(_07523_));
 sky130_fd_sc_hd__o311a_1 _28405_ (.A1(_07517_),
    .A2(\irq_mask[23] ),
    .A3(_07518_),
    .B1(_07523_),
    .C1(_07520_),
    .X(_01119_));
 sky130_fd_sc_hd__or2_1 _28406_ (.A(\irq_pending[24] ),
    .B(net17),
    .X(_07524_));
 sky130_fd_sc_hd__o311a_1 _28407_ (.A1(_07517_),
    .A2(\irq_mask[24] ),
    .A3(_07518_),
    .B1(_07524_),
    .C1(_07520_),
    .X(_01120_));
 sky130_fd_sc_hd__or2_1 _28408_ (.A(\irq_pending[25] ),
    .B(net18),
    .X(_07525_));
 sky130_fd_sc_hd__o311a_1 _28409_ (.A1(_07517_),
    .A2(\irq_mask[25] ),
    .A3(_07518_),
    .B1(_07525_),
    .C1(_07520_),
    .X(_01121_));
 sky130_fd_sc_hd__clkbuf_2 _28410_ (.A(_07475_),
    .X(_07526_));
 sky130_fd_sc_hd__clkbuf_2 _28411_ (.A(_07477_),
    .X(_07527_));
 sky130_fd_sc_hd__or2_1 _28412_ (.A(\irq_pending[26] ),
    .B(net19),
    .X(_07528_));
 sky130_fd_sc_hd__clkbuf_2 _28413_ (.A(_07327_),
    .X(_07529_));
 sky130_fd_sc_hd__o311a_1 _28414_ (.A1(_07526_),
    .A2(\irq_mask[26] ),
    .A3(_07527_),
    .B1(_07528_),
    .C1(_07529_),
    .X(_01122_));
 sky130_fd_sc_hd__or2_1 _28415_ (.A(\irq_pending[27] ),
    .B(net20),
    .X(_07530_));
 sky130_fd_sc_hd__o311a_1 _28416_ (.A1(_07526_),
    .A2(\irq_mask[27] ),
    .A3(_07527_),
    .B1(_07530_),
    .C1(_07529_),
    .X(_01123_));
 sky130_fd_sc_hd__or2_1 _28417_ (.A(\irq_pending[28] ),
    .B(net21),
    .X(_07531_));
 sky130_fd_sc_hd__o311a_1 _28418_ (.A1(_07526_),
    .A2(\irq_mask[28] ),
    .A3(_07527_),
    .B1(_07531_),
    .C1(_07529_),
    .X(_01124_));
 sky130_fd_sc_hd__or2_1 _28419_ (.A(\irq_pending[29] ),
    .B(net22),
    .X(_07532_));
 sky130_fd_sc_hd__o311a_1 _28420_ (.A1(_07526_),
    .A2(\irq_mask[29] ),
    .A3(_07527_),
    .B1(_07532_),
    .C1(_07529_),
    .X(_01125_));
 sky130_fd_sc_hd__or2_1 _28421_ (.A(\irq_pending[30] ),
    .B(net24),
    .X(_07533_));
 sky130_fd_sc_hd__o311a_1 _28422_ (.A1(_07526_),
    .A2(\irq_mask[30] ),
    .A3(_07527_),
    .B1(_07533_),
    .C1(_07529_),
    .X(_01126_));
 sky130_fd_sc_hd__or2_1 _28423_ (.A(\irq_pending[31] ),
    .B(net25),
    .X(_07534_));
 sky130_fd_sc_hd__o311a_1 _28424_ (.A1(_07526_),
    .A2(\irq_mask[31] ),
    .A3(_07527_),
    .B1(_07534_),
    .C1(_07529_),
    .X(_01127_));
 sky130_fd_sc_hd__clkbuf_2 _28425_ (.A(_06555_),
    .X(_07535_));
 sky130_fd_sc_hd__o21ai_1 _28426_ (.A1(instr_retirq),
    .A2(instr_jalr),
    .B1(_06182_),
    .Y(_07536_));
 sky130_fd_sc_hd__a21o_1 _28427_ (.A1(_06456_),
    .A2(_06182_),
    .B1(_08153_),
    .X(_07537_));
 sky130_fd_sc_hd__o211a_1 _28428_ (.A1(_07535_),
    .A2(_07536_),
    .B1(_07537_),
    .C1(_08494_),
    .X(_01128_));
 sky130_fd_sc_hd__nor4_1 _28429_ (.A(\cpu_state[0] ),
    .B(_08147_),
    .C(_07042_),
    .D(_08538_),
    .Y(_07538_));
 sky130_fd_sc_hd__o221a_1 _28430_ (.A1(is_sb_sh_sw),
    .A2(_08498_),
    .B1(_08539_),
    .B2(_08147_),
    .C1(_08296_),
    .X(_07539_));
 sky130_fd_sc_hd__o211a_1 _28431_ (.A1(_08513_),
    .A2(_08227_),
    .B1(_08319_),
    .C1(_07539_),
    .X(_07540_));
 sky130_fd_sc_hd__or4_2 _28432_ (.A(_08311_),
    .B(_08207_),
    .C(_08307_),
    .D(_06433_),
    .X(_07541_));
 sky130_fd_sc_hd__a21oi_1 _28433_ (.A1(_08312_),
    .A2(_08153_),
    .B1(_08538_),
    .Y(_07542_));
 sky130_fd_sc_hd__a31o_1 _28434_ (.A1(_07323_),
    .A2(_08305_),
    .A3(_06563_),
    .B1(_08312_),
    .X(_07543_));
 sky130_fd_sc_hd__nand4_1 _28435_ (.A(_07541_),
    .B(_07540_),
    .C(_07542_),
    .D(_07543_),
    .Y(_07544_));
 sky130_fd_sc_hd__o211a_1 _28436_ (.A1(_08522_),
    .A2(_07540_),
    .B1(_07544_),
    .C1(_08494_),
    .X(_07545_));
 sky130_fd_sc_hd__a31o_1 _28437_ (.A1(_08314_),
    .A2(_08534_),
    .A3(_07538_),
    .B1(_07545_),
    .X(_01129_));
 sky130_fd_sc_hd__a21o_1 _28438_ (.A1(_08151_),
    .A2(_08494_),
    .B1(_08174_),
    .X(_01130_));
 sky130_fd_sc_hd__or3_1 _28439_ (.A(_08163_),
    .B(_08182_),
    .C(\cpu_state[0] ),
    .X(_07546_));
 sky130_fd_sc_hd__and3b_1 _28440_ (.A_N(_07546_),
    .B(_06117_),
    .C(_08666_),
    .X(_07547_));
 sky130_fd_sc_hd__a22o_1 _28441_ (.A1(_08163_),
    .A2(_08494_),
    .B1(_07547_),
    .B2(_08160_),
    .X(_01131_));
 sky130_fd_sc_hd__nand2_1 _28442_ (.A(_08178_),
    .B(_09207_),
    .Y(_07548_));
 sky130_fd_sc_hd__clkbuf_2 _28443_ (.A(_07548_),
    .X(_07549_));
 sky130_fd_sc_hd__or3_1 _28444_ (.A(\timer[1] ),
    .B(\timer[0] ),
    .C(\timer[2] ),
    .X(_07550_));
 sky130_fd_sc_hd__or2_1 _28445_ (.A(\timer[3] ),
    .B(_07550_),
    .X(_07551_));
 sky130_fd_sc_hd__or3_1 _28446_ (.A(\timer[8] ),
    .B(_07481_),
    .C(_07551_),
    .X(_07552_));
 sky130_fd_sc_hd__or2_2 _28447_ (.A(\timer[9] ),
    .B(_07552_),
    .X(_07553_));
 sky130_fd_sc_hd__or4_1 _28448_ (.A(\timer[11] ),
    .B(\timer[10] ),
    .C(_07482_),
    .D(_07553_),
    .X(_07554_));
 sky130_fd_sc_hd__or2_1 _28449_ (.A(\timer[16] ),
    .B(_07554_),
    .X(_07555_));
 sky130_fd_sc_hd__or3_1 _28450_ (.A(\timer[17] ),
    .B(\timer[18] ),
    .C(_07555_),
    .X(_07556_));
 sky130_fd_sc_hd__or2_1 _28451_ (.A(\timer[19] ),
    .B(_07556_),
    .X(_07557_));
 sky130_fd_sc_hd__or3_1 _28452_ (.A(\timer[24] ),
    .B(_07480_),
    .C(_07557_),
    .X(_07558_));
 sky130_fd_sc_hd__or2_1 _28453_ (.A(\timer[25] ),
    .B(_07558_),
    .X(_07559_));
 sky130_fd_sc_hd__or3_2 _28454_ (.A(\timer[27] ),
    .B(\timer[26] ),
    .C(_07559_),
    .X(_07560_));
 sky130_fd_sc_hd__nor2_1 _28455_ (.A(_07479_),
    .B(_07560_),
    .Y(_07561_));
 sky130_fd_sc_hd__or2_1 _28456_ (.A(\timer[0] ),
    .B(_07561_),
    .X(_07562_));
 sky130_fd_sc_hd__and2_1 _28457_ (.A(_08178_),
    .B(_09745_),
    .X(_07563_));
 sky130_fd_sc_hd__a21o_1 _28458_ (.A1(_08635_),
    .A2(_07563_),
    .B1(_06200_),
    .X(_07564_));
 sky130_fd_sc_hd__a21oi_1 _28459_ (.A1(_07549_),
    .A2(_07562_),
    .B1(_07564_),
    .Y(_01132_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28460_ (.A(_07563_),
    .X(_07565_));
 sky130_fd_sc_hd__xnor2_1 _28461_ (.A(\timer[1] ),
    .B(_07562_),
    .Y(_07566_));
 sky130_fd_sc_hd__nand2_1 _28462_ (.A(_08744_),
    .B(_07565_),
    .Y(_07567_));
 sky130_fd_sc_hd__o211a_1 _28463_ (.A1(_07565_),
    .A2(_07566_),
    .B1(_07567_),
    .C1(_07328_),
    .X(_01133_));
 sky130_fd_sc_hd__clkbuf_2 _28464_ (.A(_07548_),
    .X(_07568_));
 sky130_fd_sc_hd__or2_1 _28465_ (.A(_08798_),
    .B(_07568_),
    .X(_07569_));
 sky130_fd_sc_hd__o21ai_1 _28466_ (.A1(\timer[1] ),
    .A2(\timer[0] ),
    .B1(\timer[2] ),
    .Y(_07570_));
 sky130_fd_sc_hd__or2_2 _28467_ (.A(_07563_),
    .B(_07561_),
    .X(_07571_));
 sky130_fd_sc_hd__clkbuf_2 _28468_ (.A(_07571_),
    .X(_07572_));
 sky130_fd_sc_hd__a21o_1 _28469_ (.A1(_07550_),
    .A2(_07570_),
    .B1(_07572_),
    .X(_07573_));
 sky130_fd_sc_hd__clkbuf_2 _28470_ (.A(_08520_),
    .X(_07574_));
 sky130_fd_sc_hd__a21oi_1 _28471_ (.A1(_07569_),
    .A2(_07573_),
    .B1(_07574_),
    .Y(_01134_));
 sky130_fd_sc_hd__buf_1 _28472_ (.A(_07548_),
    .X(_07575_));
 sky130_fd_sc_hd__or2_1 _28473_ (.A(_08865_),
    .B(_07575_),
    .X(_07576_));
 sky130_fd_sc_hd__clkbuf_2 _28474_ (.A(_07551_),
    .X(_07577_));
 sky130_fd_sc_hd__nand2_1 _28475_ (.A(\timer[3] ),
    .B(_07550_),
    .Y(_07578_));
 sky130_fd_sc_hd__a21o_1 _28476_ (.A1(_07577_),
    .A2(_07578_),
    .B1(_07572_),
    .X(_07579_));
 sky130_fd_sc_hd__clkbuf_2 _28477_ (.A(_07334_),
    .X(_07580_));
 sky130_fd_sc_hd__a21oi_1 _28478_ (.A1(_07576_),
    .A2(_07579_),
    .B1(_07580_),
    .Y(_01135_));
 sky130_fd_sc_hd__clkbuf_2 _28479_ (.A(_07571_),
    .X(_07581_));
 sky130_fd_sc_hd__nor2_1 _28480_ (.A(\timer[4] ),
    .B(_07577_),
    .Y(_07582_));
 sky130_fd_sc_hd__and2_1 _28481_ (.A(\timer[4] ),
    .B(_07577_),
    .X(_07583_));
 sky130_fd_sc_hd__nor2_1 _28482_ (.A(_07582_),
    .B(_07583_),
    .Y(_07584_));
 sky130_fd_sc_hd__o22a_1 _28483_ (.A1(_08934_),
    .A2(_07549_),
    .B1(_07581_),
    .B2(_07584_),
    .X(_07585_));
 sky130_fd_sc_hd__nor2_1 _28484_ (.A(_08521_),
    .B(_07585_),
    .Y(_01136_));
 sky130_fd_sc_hd__xnor2_1 _28485_ (.A(\timer[5] ),
    .B(_07582_),
    .Y(_07586_));
 sky130_fd_sc_hd__o22a_1 _28486_ (.A1(_08978_),
    .A2(_07549_),
    .B1(_07581_),
    .B2(_07586_),
    .X(_07587_));
 sky130_fd_sc_hd__nor2_1 _28487_ (.A(_08521_),
    .B(_07587_),
    .Y(_01137_));
 sky130_fd_sc_hd__or4_1 _28488_ (.A(\timer[5] ),
    .B(\timer[4] ),
    .C(\timer[6] ),
    .D(_07551_),
    .X(_07588_));
 sky130_fd_sc_hd__o31ai_1 _28489_ (.A1(\timer[5] ),
    .A2(\timer[4] ),
    .A3(_07577_),
    .B1(\timer[6] ),
    .Y(_07589_));
 sky130_fd_sc_hd__and2_1 _28490_ (.A(_07588_),
    .B(_07589_),
    .X(_07590_));
 sky130_fd_sc_hd__o22a_1 _28491_ (.A1(_09033_),
    .A2(_07549_),
    .B1(_07581_),
    .B2(_07590_),
    .X(_07591_));
 sky130_fd_sc_hd__nor2_1 _28492_ (.A(_08521_),
    .B(_07591_),
    .Y(_01138_));
 sky130_fd_sc_hd__clkbuf_2 _28493_ (.A(_08520_),
    .X(_07592_));
 sky130_fd_sc_hd__buf_1 _28494_ (.A(_07548_),
    .X(_07593_));
 sky130_fd_sc_hd__clkbuf_2 _28495_ (.A(_07593_),
    .X(_07594_));
 sky130_fd_sc_hd__nand2_1 _28496_ (.A(\timer[7] ),
    .B(_07588_),
    .Y(_07595_));
 sky130_fd_sc_hd__o21a_1 _28497_ (.A1(_07481_),
    .A2(_07577_),
    .B1(_07595_),
    .X(_07596_));
 sky130_fd_sc_hd__o22a_1 _28498_ (.A1(_09093_),
    .A2(_07594_),
    .B1(_07581_),
    .B2(_07596_),
    .X(_07597_));
 sky130_fd_sc_hd__nor2_1 _28499_ (.A(_07592_),
    .B(_07597_),
    .Y(_01139_));
 sky130_fd_sc_hd__or2_1 _28500_ (.A(_09151_),
    .B(_07575_),
    .X(_07598_));
 sky130_fd_sc_hd__o21ai_1 _28501_ (.A1(_07481_),
    .A2(_07577_),
    .B1(\timer[8] ),
    .Y(_07599_));
 sky130_fd_sc_hd__a21o_1 _28502_ (.A1(_07552_),
    .A2(_07599_),
    .B1(_07572_),
    .X(_07600_));
 sky130_fd_sc_hd__a21oi_1 _28503_ (.A1(_07598_),
    .A2(_07600_),
    .B1(_07580_),
    .Y(_01140_));
 sky130_fd_sc_hd__nand2_1 _28504_ (.A(\timer[9] ),
    .B(_07552_),
    .Y(_07601_));
 sky130_fd_sc_hd__clkbuf_2 _28505_ (.A(_07571_),
    .X(_07602_));
 sky130_fd_sc_hd__a21o_1 _28506_ (.A1(_07553_),
    .A2(_07601_),
    .B1(_07602_),
    .X(_07603_));
 sky130_fd_sc_hd__or2_1 _28507_ (.A(_09205_),
    .B(_07575_),
    .X(_07604_));
 sky130_fd_sc_hd__a21oi_1 _28508_ (.A1(_07603_),
    .A2(_07604_),
    .B1(_07580_),
    .Y(_01141_));
 sky130_fd_sc_hd__xor2_1 _28509_ (.A(_09247_),
    .B(_07553_),
    .X(_07605_));
 sky130_fd_sc_hd__o22a_1 _28510_ (.A1(_09245_),
    .A2(_07594_),
    .B1(_07581_),
    .B2(_07605_),
    .X(_07606_));
 sky130_fd_sc_hd__nor2_1 _28511_ (.A(_07592_),
    .B(_07606_),
    .Y(_01142_));
 sky130_fd_sc_hd__nor3_1 _28512_ (.A(\timer[11] ),
    .B(_09247_),
    .C(_07553_),
    .Y(_07607_));
 sky130_fd_sc_hd__o21a_1 _28513_ (.A1(_09247_),
    .A2(_07553_),
    .B1(\timer[11] ),
    .X(_07608_));
 sky130_fd_sc_hd__nor2_1 _28514_ (.A(_07607_),
    .B(_07608_),
    .Y(_07609_));
 sky130_fd_sc_hd__o22a_1 _28515_ (.A1(_09282_),
    .A2(_07594_),
    .B1(_07581_),
    .B2(_07609_),
    .X(_07610_));
 sky130_fd_sc_hd__nor2_1 _28516_ (.A(_07592_),
    .B(_07610_),
    .Y(_01143_));
 sky130_fd_sc_hd__clkbuf_2 _28517_ (.A(_07571_),
    .X(_07611_));
 sky130_fd_sc_hd__xnor2_1 _28518_ (.A(\timer[12] ),
    .B(_07607_),
    .Y(_07612_));
 sky130_fd_sc_hd__o22a_1 _28519_ (.A1(_09332_),
    .A2(_07594_),
    .B1(_07611_),
    .B2(_07612_),
    .X(_07613_));
 sky130_fd_sc_hd__nor2_1 _28520_ (.A(_07592_),
    .B(_07613_),
    .Y(_01144_));
 sky130_fd_sc_hd__or4_1 _28521_ (.A(\timer[11] ),
    .B(_09247_),
    .C(\timer[12] ),
    .D(_07553_),
    .X(_07614_));
 sky130_fd_sc_hd__nor2_1 _28522_ (.A(\timer[13] ),
    .B(_07614_),
    .Y(_07615_));
 sky130_fd_sc_hd__and2_1 _28523_ (.A(\timer[13] ),
    .B(_07614_),
    .X(_07616_));
 sky130_fd_sc_hd__nor2_1 _28524_ (.A(_07615_),
    .B(_07616_),
    .Y(_07617_));
 sky130_fd_sc_hd__o22a_1 _28525_ (.A1(_09372_),
    .A2(_07594_),
    .B1(_07611_),
    .B2(_07617_),
    .X(_07618_));
 sky130_fd_sc_hd__nor2_1 _28526_ (.A(_07592_),
    .B(_07618_),
    .Y(_01145_));
 sky130_fd_sc_hd__xnor2_1 _28527_ (.A(\timer[14] ),
    .B(_07615_),
    .Y(_07619_));
 sky130_fd_sc_hd__o22a_1 _28528_ (.A1(_09414_),
    .A2(_07594_),
    .B1(_07611_),
    .B2(_07619_),
    .X(_07620_));
 sky130_fd_sc_hd__nor2_1 _28529_ (.A(_07592_),
    .B(_07620_),
    .Y(_01146_));
 sky130_fd_sc_hd__o31ai_1 _28530_ (.A1(\timer[13] ),
    .A2(\timer[14] ),
    .A3(_07614_),
    .B1(\timer[15] ),
    .Y(_07621_));
 sky130_fd_sc_hd__a21o_1 _28531_ (.A1(_07554_),
    .A2(_07621_),
    .B1(_07602_),
    .X(_07622_));
 sky130_fd_sc_hd__or2_1 _28532_ (.A(_09453_),
    .B(_07575_),
    .X(_07623_));
 sky130_fd_sc_hd__a21oi_1 _28533_ (.A1(_07622_),
    .A2(_07623_),
    .B1(_07580_),
    .Y(_01147_));
 sky130_fd_sc_hd__nand2_1 _28534_ (.A(\timer[16] ),
    .B(_07554_),
    .Y(_07624_));
 sky130_fd_sc_hd__a21o_1 _28535_ (.A1(_07555_),
    .A2(_07624_),
    .B1(_07602_),
    .X(_07625_));
 sky130_fd_sc_hd__or2_1 _28536_ (.A(_09507_),
    .B(_07575_),
    .X(_07626_));
 sky130_fd_sc_hd__a21oi_1 _28537_ (.A1(_07625_),
    .A2(_07626_),
    .B1(_07580_),
    .Y(_01148_));
 sky130_fd_sc_hd__xor2_1 _28538_ (.A(\timer[17] ),
    .B(_07555_),
    .X(_07627_));
 sky130_fd_sc_hd__o22a_1 _28539_ (.A1(_09545_),
    .A2(_07568_),
    .B1(_07611_),
    .B2(_07627_),
    .X(_07628_));
 sky130_fd_sc_hd__nor2_1 _28540_ (.A(_07574_),
    .B(_07628_),
    .Y(_01149_));
 sky130_fd_sc_hd__o21ai_1 _28541_ (.A1(\timer[17] ),
    .A2(_07555_),
    .B1(\timer[18] ),
    .Y(_07629_));
 sky130_fd_sc_hd__a21o_1 _28542_ (.A1(_07556_),
    .A2(_07629_),
    .B1(_07602_),
    .X(_07630_));
 sky130_fd_sc_hd__or2_1 _28543_ (.A(_09589_),
    .B(_07575_),
    .X(_07631_));
 sky130_fd_sc_hd__a21oi_1 _28544_ (.A1(_07630_),
    .A2(_07631_),
    .B1(_07580_),
    .Y(_01150_));
 sky130_fd_sc_hd__clkbuf_2 _28545_ (.A(_07557_),
    .X(_07632_));
 sky130_fd_sc_hd__nand2_1 _28546_ (.A(\timer[19] ),
    .B(_07556_),
    .Y(_07633_));
 sky130_fd_sc_hd__a21o_1 _28547_ (.A1(_07632_),
    .A2(_07633_),
    .B1(_07602_),
    .X(_07634_));
 sky130_fd_sc_hd__or2_1 _28548_ (.A(_09626_),
    .B(_07593_),
    .X(_07635_));
 sky130_fd_sc_hd__a21oi_1 _28549_ (.A1(_07634_),
    .A2(_07635_),
    .B1(_07335_),
    .Y(_01151_));
 sky130_fd_sc_hd__xor2_1 _28550_ (.A(\timer[20] ),
    .B(_07632_),
    .X(_07636_));
 sky130_fd_sc_hd__o22a_1 _28551_ (.A1(_09667_),
    .A2(_07568_),
    .B1(_07611_),
    .B2(_07636_),
    .X(_07637_));
 sky130_fd_sc_hd__nor2_1 _28552_ (.A(_07574_),
    .B(_07637_),
    .Y(_01152_));
 sky130_fd_sc_hd__or3_1 _28553_ (.A(\timer[21] ),
    .B(\timer[20] ),
    .C(_07632_),
    .X(_07638_));
 sky130_fd_sc_hd__o21ai_1 _28554_ (.A1(\timer[20] ),
    .A2(_07632_),
    .B1(\timer[21] ),
    .Y(_07639_));
 sky130_fd_sc_hd__a21o_1 _28555_ (.A1(_07638_),
    .A2(_07639_),
    .B1(_07602_),
    .X(_07640_));
 sky130_fd_sc_hd__or2_1 _28556_ (.A(_09704_),
    .B(_07593_),
    .X(_07641_));
 sky130_fd_sc_hd__a21oi_1 _28557_ (.A1(_07640_),
    .A2(_07641_),
    .B1(_07335_),
    .Y(_01153_));
 sky130_fd_sc_hd__xor2_1 _28558_ (.A(\timer[22] ),
    .B(_07638_),
    .X(_07642_));
 sky130_fd_sc_hd__o22a_1 _28559_ (.A1(_09744_),
    .A2(_07568_),
    .B1(_07611_),
    .B2(_07642_),
    .X(_07643_));
 sky130_fd_sc_hd__nor2_1 _28560_ (.A(_07574_),
    .B(_07643_),
    .Y(_01154_));
 sky130_fd_sc_hd__o21ai_1 _28561_ (.A1(\timer[22] ),
    .A2(_07638_),
    .B1(\timer[23] ),
    .Y(_07644_));
 sky130_fd_sc_hd__o21a_1 _28562_ (.A1(_07480_),
    .A2(_07632_),
    .B1(_07644_),
    .X(_07645_));
 sky130_fd_sc_hd__o22a_1 _28563_ (.A1(_09781_),
    .A2(_07568_),
    .B1(_07571_),
    .B2(_07645_),
    .X(_07646_));
 sky130_fd_sc_hd__nor2_1 _28564_ (.A(_07574_),
    .B(_07646_),
    .Y(_01155_));
 sky130_fd_sc_hd__o21ai_1 _28565_ (.A1(_07480_),
    .A2(_07632_),
    .B1(\timer[24] ),
    .Y(_07647_));
 sky130_fd_sc_hd__a21o_1 _28566_ (.A1(_07558_),
    .A2(_07647_),
    .B1(_07572_),
    .X(_07648_));
 sky130_fd_sc_hd__or2_1 _28567_ (.A(_09821_),
    .B(_07593_),
    .X(_07649_));
 sky130_fd_sc_hd__a21oi_1 _28568_ (.A1(_07648_),
    .A2(_07649_),
    .B1(_07335_),
    .Y(_01156_));
 sky130_fd_sc_hd__nand2_1 _28569_ (.A(\timer[25] ),
    .B(_07558_),
    .Y(_07650_));
 sky130_fd_sc_hd__a21o_1 _28570_ (.A1(_07559_),
    .A2(_07650_),
    .B1(_07572_),
    .X(_07651_));
 sky130_fd_sc_hd__or2_1 _28571_ (.A(_09855_),
    .B(_07593_),
    .X(_07652_));
 sky130_fd_sc_hd__a21oi_1 _28572_ (.A1(_07651_),
    .A2(_07652_),
    .B1(_07335_),
    .Y(_01157_));
 sky130_fd_sc_hd__xor2_1 _28573_ (.A(\timer[26] ),
    .B(_07559_),
    .X(_07653_));
 sky130_fd_sc_hd__o22a_1 _28574_ (.A1(_09888_),
    .A2(_07568_),
    .B1(_07571_),
    .B2(_07653_),
    .X(_07654_));
 sky130_fd_sc_hd__nor2_1 _28575_ (.A(_07574_),
    .B(_07654_),
    .Y(_01158_));
 sky130_fd_sc_hd__and2b_1 _28576_ (.A_N(_07560_),
    .B(_07479_),
    .X(_07655_));
 sky130_fd_sc_hd__o21a_1 _28577_ (.A1(\timer[26] ),
    .A2(_07559_),
    .B1(\timer[27] ),
    .X(_07656_));
 sky130_fd_sc_hd__nand2_1 _28578_ (.A(_09929_),
    .B(_07565_),
    .Y(_07657_));
 sky130_fd_sc_hd__o311a_1 _28579_ (.A1(_07565_),
    .A2(_07655_),
    .A3(_07656_),
    .B1(_07657_),
    .C1(_06184_),
    .X(_01159_));
 sky130_fd_sc_hd__xnor2_1 _28580_ (.A(\timer[28] ),
    .B(_07560_),
    .Y(_07658_));
 sky130_fd_sc_hd__a21o_1 _28581_ (.A1(_07479_),
    .A2(_07658_),
    .B1(_07563_),
    .X(_07659_));
 sky130_fd_sc_hd__o211a_1 _28582_ (.A1(_07467_),
    .A2(_07549_),
    .B1(_07659_),
    .C1(_07328_),
    .X(_01160_));
 sky130_fd_sc_hd__or3_1 _28583_ (.A(\timer[29] ),
    .B(\timer[28] ),
    .C(_07560_),
    .X(_07660_));
 sky130_fd_sc_hd__o21ba_1 _28584_ (.A1(\timer[31] ),
    .A2(\timer[30] ),
    .B1_N(_07660_),
    .X(_07661_));
 sky130_fd_sc_hd__o21a_1 _28585_ (.A1(\timer[28] ),
    .A2(_07560_),
    .B1(\timer[29] ),
    .X(_07662_));
 sky130_fd_sc_hd__nand2_1 _28586_ (.A(_10003_),
    .B(_07565_),
    .Y(_07663_));
 sky130_fd_sc_hd__o311a_1 _28587_ (.A1(_07565_),
    .A2(_07661_),
    .A3(_07662_),
    .B1(_07663_),
    .C1(_06184_),
    .X(_01161_));
 sky130_fd_sc_hd__or2_1 _28588_ (.A(\timer[30] ),
    .B(_07660_),
    .X(_07664_));
 sky130_fd_sc_hd__nand2_1 _28589_ (.A(\timer[30] ),
    .B(_07660_),
    .Y(_07665_));
 sky130_fd_sc_hd__a21o_1 _28590_ (.A1(_07664_),
    .A2(_07665_),
    .B1(_07572_),
    .X(_07666_));
 sky130_fd_sc_hd__or2_1 _28591_ (.A(_10040_),
    .B(_07593_),
    .X(_07667_));
 sky130_fd_sc_hd__a21oi_1 _28592_ (.A1(_07666_),
    .A2(_07667_),
    .B1(_07335_),
    .Y(_01162_));
 sky130_fd_sc_hd__a21o_1 _28593_ (.A1(\timer[31] ),
    .A2(_07664_),
    .B1(_07563_),
    .X(_07668_));
 sky130_fd_sc_hd__o211a_1 _28594_ (.A1(_07473_),
    .A2(_07549_),
    .B1(_07668_),
    .C1(_07328_),
    .X(_01163_));
 sky130_fd_sc_hd__nor2_1 _28595_ (.A(_10305_),
    .B(_05052_),
    .Y(_07669_));
 sky130_fd_sc_hd__a32o_1 _28596_ (.A1(_06333_),
    .A2(_08277_),
    .A3(_07669_),
    .B1(_06346_),
    .B2(_05052_),
    .X(_01164_));
 sky130_fd_sc_hd__xor2_1 _28597_ (.A(_10305_),
    .B(_08232_),
    .X(_07670_));
 sky130_fd_sc_hd__and3_1 _28598_ (.A(_06129_),
    .B(_07324_),
    .C(_07670_),
    .X(_07671_));
 sky130_fd_sc_hd__clkbuf_1 _28599_ (.A(_07671_),
    .X(_01165_));
 sky130_fd_sc_hd__o211a_1 _28600_ (.A1(\cpu_state[1] ),
    .A2(_08540_),
    .B1(_08514_),
    .C1(_08495_),
    .X(_07672_));
 sky130_fd_sc_hd__and3_1 _28601_ (.A(_08319_),
    .B(_08498_),
    .C(_07672_),
    .X(_07673_));
 sky130_fd_sc_hd__o21a_1 _28602_ (.A1(_08313_),
    .A2(_08534_),
    .B1(_08311_),
    .X(_07674_));
 sky130_fd_sc_hd__a211o_1 _28603_ (.A1(_08295_),
    .A2(_06451_),
    .B1(_08538_),
    .C1(_08671_),
    .X(_07675_));
 sky130_fd_sc_hd__or3b_1 _28604_ (.A(_07674_),
    .B(_07675_),
    .C_N(_07673_),
    .X(_07676_));
 sky130_fd_sc_hd__o211a_1 _28605_ (.A1(_10317_),
    .A2(_07673_),
    .B1(_07676_),
    .C1(_07328_),
    .X(_01166_));
 sky130_fd_sc_hd__o21a_1 _28606_ (.A1(_08873_),
    .A2(_06117_),
    .B1(_04984_),
    .X(_07677_));
 sky130_fd_sc_hd__o21a_1 _28607_ (.A1(_08297_),
    .A2(_07677_),
    .B1(_06130_),
    .X(_01167_));
 sky130_fd_sc_hd__o21ai_1 _28608_ (.A1(_08294_),
    .A2(instr_jalr),
    .B1(_07674_),
    .Y(_07678_));
 sky130_fd_sc_hd__or2_1 _28609_ (.A(_08311_),
    .B(_06118_),
    .X(_07679_));
 sky130_fd_sc_hd__and4_1 _28610_ (.A(_06124_),
    .B(_08495_),
    .C(_07678_),
    .D(_07679_),
    .X(_07680_));
 sky130_fd_sc_hd__nand2_1 _28611_ (.A(_07541_),
    .B(_07680_),
    .Y(_07681_));
 sky130_fd_sc_hd__a31o_1 _28612_ (.A1(_08495_),
    .A2(_06119_),
    .A3(_07679_),
    .B1(_10316_),
    .X(_07682_));
 sky130_fd_sc_hd__and3_1 _28613_ (.A(_06129_),
    .B(_07681_),
    .C(_07682_),
    .X(_07683_));
 sky130_fd_sc_hd__clkbuf_1 _28614_ (.A(_07683_),
    .X(_01168_));
 sky130_fd_sc_hd__nor2_1 _28615_ (.A(_08232_),
    .B(_09048_),
    .Y(_07684_));
 sky130_fd_sc_hd__o21a_1 _28616_ (.A1(_08168_),
    .A2(_07684_),
    .B1(_08322_),
    .X(_07685_));
 sky130_fd_sc_hd__a22o_1 _28617_ (.A1(instr_lh),
    .A2(_08174_),
    .B1(_07685_),
    .B2(latched_is_lh),
    .X(_01170_));
 sky130_fd_sc_hd__a22o_1 _28618_ (.A1(instr_lb),
    .A2(_08174_),
    .B1(_07685_),
    .B2(latched_is_lb),
    .X(_01171_));
 sky130_fd_sc_hd__or3_1 _28619_ (.A(\pcpi_timeout_counter[2] ),
    .B(\pcpi_timeout_counter[1] ),
    .C(\pcpi_timeout_counter[0] ),
    .X(_07686_));
 sky130_fd_sc_hd__nor2_1 _28620_ (.A(\pcpi_timeout_counter[3] ),
    .B(_07686_),
    .Y(_07687_));
 sky130_fd_sc_hd__o21bai_1 _28621_ (.A1(\pcpi_timeout_counter[0] ),
    .A2(_07687_),
    .B1_N(_08137_),
    .Y(_01172_));
 sky130_fd_sc_hd__nor3_1 _28622_ (.A(\pcpi_timeout_counter[1] ),
    .B(\pcpi_timeout_counter[0] ),
    .C(_07687_),
    .Y(_07688_));
 sky130_fd_sc_hd__a211o_1 _28623_ (.A1(\pcpi_timeout_counter[1] ),
    .A2(\pcpi_timeout_counter[0] ),
    .B1(_08137_),
    .C1(_07688_),
    .X(_01173_));
 sky130_vsdinv _28624_ (.A(_07686_),
    .Y(_07689_));
 sky130_fd_sc_hd__o21a_1 _28625_ (.A1(\pcpi_timeout_counter[1] ),
    .A2(\pcpi_timeout_counter[0] ),
    .B1(\pcpi_timeout_counter[2] ),
    .X(_07690_));
 sky130_fd_sc_hd__a211o_1 _28626_ (.A1(net466),
    .A2(_07689_),
    .B1(_07690_),
    .C1(_08137_),
    .X(_01174_));
 sky130_fd_sc_hd__a21o_1 _28627_ (.A1(net466),
    .A2(_07686_),
    .B1(_08137_),
    .X(_01175_));
 sky130_fd_sc_hd__and2_1 _28628_ (.A(_06114_),
    .B(_07687_),
    .X(_07691_));
 sky130_fd_sc_hd__clkbuf_1 _28629_ (.A(_07691_),
    .X(_01176_));
 sky130_fd_sc_hd__and4b_1 _28630_ (.A_N(_08277_),
    .B(_07669_),
    .C(_06532_),
    .D(_08176_),
    .X(_07692_));
 sky130_fd_sc_hd__clkbuf_1 _28631_ (.A(_07692_),
    .X(_01177_));
 sky130_fd_sc_hd__nor2_2 _28632_ (.A(_06473_),
    .B(decoder_pseudo_trigger),
    .Y(_07693_));
 sky130_fd_sc_hd__buf_2 _28633_ (.A(_07693_),
    .X(_07694_));
 sky130_fd_sc_hd__buf_2 _28634_ (.A(_07694_),
    .X(_07695_));
 sky130_fd_sc_hd__mux2_1 _28635_ (.A0(net235),
    .A1(\mem_rdata_q[0] ),
    .S(_07695_),
    .X(_07696_));
 sky130_fd_sc_hd__clkbuf_1 _28636_ (.A(_07696_),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_1 _28637_ (.A0(net246),
    .A1(\mem_rdata_q[1] ),
    .S(_07695_),
    .X(_07697_));
 sky130_fd_sc_hd__clkbuf_1 _28638_ (.A(_07697_),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_1 _28639_ (.A0(net257),
    .A1(\mem_rdata_q[2] ),
    .S(_07695_),
    .X(_07698_));
 sky130_fd_sc_hd__clkbuf_1 _28640_ (.A(_07698_),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _28641_ (.A0(net260),
    .A1(\mem_rdata_q[3] ),
    .S(_07695_),
    .X(_07699_));
 sky130_fd_sc_hd__clkbuf_1 _28642_ (.A(_07699_),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _28643_ (.A0(net261),
    .A1(\mem_rdata_q[4] ),
    .S(_07695_),
    .X(_07700_));
 sky130_fd_sc_hd__clkbuf_1 _28644_ (.A(_07700_),
    .X(_01182_));
 sky130_fd_sc_hd__clkbuf_2 _28645_ (.A(_07693_),
    .X(_07701_));
 sky130_fd_sc_hd__clkbuf_4 _28646_ (.A(_07701_),
    .X(_07702_));
 sky130_fd_sc_hd__mux2_1 _28647_ (.A0(net262),
    .A1(\mem_rdata_q[5] ),
    .S(_07702_),
    .X(_07703_));
 sky130_fd_sc_hd__clkbuf_1 _28648_ (.A(_07703_),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _28649_ (.A0(net263),
    .A1(\mem_rdata_q[6] ),
    .S(_07702_),
    .X(_07704_));
 sky130_fd_sc_hd__clkbuf_1 _28650_ (.A(_07704_),
    .X(_01184_));
 sky130_fd_sc_hd__or2_4 _28651_ (.A(_08233_),
    .B(decoder_pseudo_trigger),
    .X(_07705_));
 sky130_fd_sc_hd__clkbuf_2 _28652_ (.A(_07705_),
    .X(_07706_));
 sky130_fd_sc_hd__mux2_1 _28653_ (.A0(\mem_rdata_q[7] ),
    .A1(net264),
    .S(_07706_),
    .X(_07707_));
 sky130_fd_sc_hd__clkbuf_1 _28654_ (.A(_07707_),
    .X(_01185_));
 sky130_fd_sc_hd__clkbuf_2 _28655_ (.A(_07705_),
    .X(_07708_));
 sky130_fd_sc_hd__mux2_1 _28656_ (.A0(\mem_rdata_q[8] ),
    .A1(net265),
    .S(_07708_),
    .X(_07709_));
 sky130_fd_sc_hd__clkbuf_1 _28657_ (.A(_07709_),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _28658_ (.A0(\mem_rdata_q[9] ),
    .A1(net266),
    .S(_07708_),
    .X(_07710_));
 sky130_fd_sc_hd__clkbuf_1 _28659_ (.A(_07710_),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _28660_ (.A0(\mem_rdata_q[10] ),
    .A1(net236),
    .S(_07708_),
    .X(_07711_));
 sky130_fd_sc_hd__clkbuf_1 _28661_ (.A(_07711_),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _28662_ (.A0(\mem_rdata_q[11] ),
    .A1(net237),
    .S(_07708_),
    .X(_07712_));
 sky130_fd_sc_hd__clkbuf_1 _28663_ (.A(_07712_),
    .X(_01189_));
 sky130_fd_sc_hd__buf_2 _28664_ (.A(\mem_rdata_q[12] ),
    .X(_07713_));
 sky130_fd_sc_hd__mux2_1 _28665_ (.A0(net238),
    .A1(_07713_),
    .S(_07702_),
    .X(_07714_));
 sky130_fd_sc_hd__clkbuf_1 _28666_ (.A(_07714_),
    .X(_01190_));
 sky130_fd_sc_hd__buf_2 _28667_ (.A(\mem_rdata_q[13] ),
    .X(_07715_));
 sky130_fd_sc_hd__mux2_1 _28668_ (.A0(net239),
    .A1(_07715_),
    .S(_07702_),
    .X(_07716_));
 sky130_fd_sc_hd__clkbuf_1 _28669_ (.A(_07716_),
    .X(_01191_));
 sky130_fd_sc_hd__buf_2 _28670_ (.A(\mem_rdata_q[14] ),
    .X(_07717_));
 sky130_fd_sc_hd__mux2_1 _28671_ (.A0(net240),
    .A1(_07717_),
    .S(_07702_),
    .X(_07718_));
 sky130_fd_sc_hd__clkbuf_1 _28672_ (.A(_07718_),
    .X(_01192_));
 sky130_fd_sc_hd__mux2_1 _28673_ (.A0(\mem_rdata_q[15] ),
    .A1(net241),
    .S(_07708_),
    .X(_07719_));
 sky130_fd_sc_hd__clkbuf_1 _28674_ (.A(_07719_),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_1 _28675_ (.A0(\mem_rdata_q[16] ),
    .A1(net242),
    .S(_07708_),
    .X(_07720_));
 sky130_fd_sc_hd__clkbuf_1 _28676_ (.A(_07720_),
    .X(_01194_));
 sky130_fd_sc_hd__clkbuf_2 _28677_ (.A(_07705_),
    .X(_07721_));
 sky130_fd_sc_hd__mux2_1 _28678_ (.A0(\mem_rdata_q[17] ),
    .A1(net243),
    .S(_07721_),
    .X(_07722_));
 sky130_fd_sc_hd__clkbuf_1 _28679_ (.A(_07722_),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_1 _28680_ (.A0(\mem_rdata_q[18] ),
    .A1(net244),
    .S(_07721_),
    .X(_07723_));
 sky130_fd_sc_hd__clkbuf_1 _28681_ (.A(_07723_),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_1 _28682_ (.A0(\mem_rdata_q[19] ),
    .A1(net245),
    .S(_07721_),
    .X(_07724_));
 sky130_fd_sc_hd__clkbuf_1 _28683_ (.A(_07724_),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _28684_ (.A0(\mem_rdata_q[20] ),
    .A1(net247),
    .S(_07721_),
    .X(_07725_));
 sky130_fd_sc_hd__clkbuf_1 _28685_ (.A(_07725_),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_1 _28686_ (.A0(\mem_rdata_q[21] ),
    .A1(net248),
    .S(_07721_),
    .X(_07726_));
 sky130_fd_sc_hd__clkbuf_1 _28687_ (.A(_07726_),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_1 _28688_ (.A0(\mem_rdata_q[22] ),
    .A1(net249),
    .S(_07721_),
    .X(_07727_));
 sky130_fd_sc_hd__clkbuf_1 _28689_ (.A(_07727_),
    .X(_01200_));
 sky130_fd_sc_hd__clkbuf_2 _28690_ (.A(_07705_),
    .X(_07728_));
 sky130_fd_sc_hd__buf_2 _28691_ (.A(_07728_),
    .X(_07729_));
 sky130_fd_sc_hd__mux2_1 _28692_ (.A0(\mem_rdata_q[23] ),
    .A1(net250),
    .S(_07729_),
    .X(_07730_));
 sky130_fd_sc_hd__clkbuf_1 _28693_ (.A(_07730_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _28694_ (.A0(\mem_rdata_q[24] ),
    .A1(net251),
    .S(_07729_),
    .X(_07731_));
 sky130_fd_sc_hd__clkbuf_1 _28695_ (.A(_07731_),
    .X(_01202_));
 sky130_fd_sc_hd__clkbuf_2 _28696_ (.A(\mem_rdata_q[25] ),
    .X(_07732_));
 sky130_fd_sc_hd__mux2_1 _28697_ (.A0(net252),
    .A1(_07732_),
    .S(_07702_),
    .X(_07733_));
 sky130_fd_sc_hd__clkbuf_1 _28698_ (.A(_07733_),
    .X(_01203_));
 sky130_fd_sc_hd__clkbuf_2 _28699_ (.A(\mem_rdata_q[26] ),
    .X(_07734_));
 sky130_fd_sc_hd__mux2_1 _28700_ (.A0(_07734_),
    .A1(net253),
    .S(_07729_),
    .X(_07735_));
 sky130_fd_sc_hd__clkbuf_1 _28701_ (.A(_07735_),
    .X(_01204_));
 sky130_fd_sc_hd__buf_2 _28702_ (.A(\mem_rdata_q[27] ),
    .X(_07736_));
 sky130_fd_sc_hd__mux2_1 _28703_ (.A0(_07736_),
    .A1(net254),
    .S(_07729_),
    .X(_07737_));
 sky130_fd_sc_hd__clkbuf_1 _28704_ (.A(_07737_),
    .X(_01205_));
 sky130_fd_sc_hd__buf_1 _28705_ (.A(_07701_),
    .X(_07738_));
 sky130_fd_sc_hd__clkbuf_2 _28706_ (.A(_07738_),
    .X(_07739_));
 sky130_fd_sc_hd__buf_2 _28707_ (.A(_07739_),
    .X(_07740_));
 sky130_fd_sc_hd__nor2_1 _28708_ (.A(\mem_rdata_q[28] ),
    .B(_07728_),
    .Y(_07741_));
 sky130_fd_sc_hd__o21ba_1 _28709_ (.A1(net255),
    .A2(_07740_),
    .B1_N(_07741_),
    .X(_01206_));
 sky130_fd_sc_hd__clkbuf_2 _28710_ (.A(\mem_rdata_q[29] ),
    .X(_07742_));
 sky130_fd_sc_hd__buf_2 _28711_ (.A(_07694_),
    .X(_07743_));
 sky130_fd_sc_hd__mux2_1 _28712_ (.A0(net256),
    .A1(_07742_),
    .S(_07743_),
    .X(_07744_));
 sky130_fd_sc_hd__clkbuf_1 _28713_ (.A(_07744_),
    .X(_01207_));
 sky130_fd_sc_hd__clkbuf_2 _28714_ (.A(\mem_rdata_q[30] ),
    .X(_07745_));
 sky130_fd_sc_hd__mux2_1 _28715_ (.A0(net258),
    .A1(_07745_),
    .S(_07743_),
    .X(_07746_));
 sky130_fd_sc_hd__clkbuf_1 _28716_ (.A(_07746_),
    .X(_01208_));
 sky130_fd_sc_hd__clkbuf_2 _28717_ (.A(\mem_rdata_q[31] ),
    .X(_07747_));
 sky130_fd_sc_hd__mux2_1 _28718_ (.A0(net259),
    .A1(_07747_),
    .S(_07743_),
    .X(_07748_));
 sky130_fd_sc_hd__clkbuf_1 _28719_ (.A(_07748_),
    .X(_01209_));
 sky130_fd_sc_hd__buf_2 _28720_ (.A(_08535_),
    .X(_07749_));
 sky130_fd_sc_hd__and3_1 _28721_ (.A(_00613_),
    .B(_00614_),
    .C(_00615_),
    .X(_07750_));
 sky130_fd_sc_hd__and2b_1 _28722_ (.A_N(_00616_),
    .B(_07750_),
    .X(_07751_));
 sky130_fd_sc_hd__nor2_1 _28723_ (.A(_08535_),
    .B(_00619_),
    .Y(_07752_));
 sky130_fd_sc_hd__and3_1 _28724_ (.A(_00617_),
    .B(_00618_),
    .C(_07752_),
    .X(_07753_));
 sky130_fd_sc_hd__a22o_1 _28725_ (.A1(instr_lui),
    .A2(_07749_),
    .B1(_07751_),
    .B2(_07753_),
    .X(_01210_));
 sky130_fd_sc_hd__and3b_1 _28726_ (.A_N(_00618_),
    .B(_07752_),
    .C(_00617_),
    .X(_07754_));
 sky130_fd_sc_hd__a22o_1 _28727_ (.A1(instr_auipc),
    .A2(_07749_),
    .B1(_07751_),
    .B2(_07754_),
    .X(_01211_));
 sky130_fd_sc_hd__and3b_1 _28728_ (.A_N(_00617_),
    .B(_00618_),
    .C(_00619_),
    .X(_07755_));
 sky130_fd_sc_hd__and3_1 _28729_ (.A(_05537_),
    .B(_07750_),
    .C(_07755_),
    .X(_07756_));
 sky130_fd_sc_hd__a22o_1 _28730_ (.A1(_07535_),
    .A2(_07749_),
    .B1(_00616_),
    .B2(_07756_),
    .X(_01212_));
 sky130_fd_sc_hd__nor2_1 _28731_ (.A(_08182_),
    .B(_07701_),
    .Y(_07757_));
 sky130_fd_sc_hd__clkbuf_2 _28732_ (.A(_07757_),
    .X(_07758_));
 sky130_fd_sc_hd__clkbuf_2 _28733_ (.A(_07758_),
    .X(_07759_));
 sky130_fd_sc_hd__nor3_1 _28734_ (.A(\mem_rdata_q[14] ),
    .B(\mem_rdata_q[13] ),
    .C(\mem_rdata_q[12] ),
    .Y(_07760_));
 sky130_fd_sc_hd__and3_1 _28735_ (.A(_08294_),
    .B(_08321_),
    .C(_07694_),
    .X(_07761_));
 sky130_fd_sc_hd__clkbuf_2 _28736_ (.A(_07761_),
    .X(_07762_));
 sky130_fd_sc_hd__a22o_1 _28737_ (.A1(net447),
    .A2(_07759_),
    .B1(net372),
    .B2(_07762_),
    .X(_01213_));
 sky130_fd_sc_hd__or2b_1 _28738_ (.A(\mem_rdata_q[13] ),
    .B_N(\mem_rdata_q[12] ),
    .X(_07763_));
 sky130_fd_sc_hd__nor2_2 _28739_ (.A(\mem_rdata_q[14] ),
    .B(_07763_),
    .Y(_07764_));
 sky130_fd_sc_hd__a22o_1 _28740_ (.A1(instr_bne),
    .A2(_07759_),
    .B1(_07762_),
    .B2(_07764_),
    .X(_01214_));
 sky130_fd_sc_hd__nor3b_2 _28741_ (.A(_07715_),
    .B(_07713_),
    .C_N(_07717_),
    .Y(_07765_));
 sky130_fd_sc_hd__a22o_1 _28742_ (.A1(instr_blt),
    .A2(_07759_),
    .B1(_07762_),
    .B2(_07765_),
    .X(_01215_));
 sky130_fd_sc_hd__and3b_1 _28743_ (.A_N(\mem_rdata_q[13] ),
    .B(\mem_rdata_q[12] ),
    .C(\mem_rdata_q[14] ),
    .X(_07766_));
 sky130_fd_sc_hd__clkbuf_2 _28744_ (.A(_07766_),
    .X(_07767_));
 sky130_fd_sc_hd__a22o_1 _28745_ (.A1(instr_bge),
    .A2(_07759_),
    .B1(_07762_),
    .B2(_07767_),
    .X(_01216_));
 sky130_fd_sc_hd__and3b_1 _28746_ (.A_N(_07713_),
    .B(_07715_),
    .C(_07717_),
    .X(_07768_));
 sky130_fd_sc_hd__a22o_1 _28747_ (.A1(net468),
    .A2(_07759_),
    .B1(_07762_),
    .B2(_07768_),
    .X(_01217_));
 sky130_fd_sc_hd__clkbuf_2 _28748_ (.A(_07757_),
    .X(_07769_));
 sky130_fd_sc_hd__and3_1 _28749_ (.A(_07717_),
    .B(_07715_),
    .C(_07713_),
    .X(_07770_));
 sky130_fd_sc_hd__a22o_1 _28750_ (.A1(instr_bgeu),
    .A2(_07769_),
    .B1(_07762_),
    .B2(_07770_),
    .X(_01218_));
 sky130_fd_sc_hd__clkbuf_2 _28751_ (.A(_08535_),
    .X(_07771_));
 sky130_fd_sc_hd__or4b_1 _28752_ (.A(_00625_),
    .B(_00626_),
    .C(_00627_),
    .D_N(_07755_),
    .X(_07772_));
 sky130_fd_sc_hd__nor2_1 _28753_ (.A(_08536_),
    .B(_07772_),
    .Y(_07773_));
 sky130_fd_sc_hd__a22o_1 _28754_ (.A1(instr_jalr),
    .A2(_07771_),
    .B1(_07751_),
    .B2(_07773_),
    .X(_01219_));
 sky130_fd_sc_hd__clkbuf_2 _28755_ (.A(_07706_),
    .X(_07774_));
 sky130_fd_sc_hd__and2_1 _28756_ (.A(is_lb_lh_lw_lbu_lhu),
    .B(_07694_),
    .X(_07775_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28757_ (.A(_07775_),
    .X(_07776_));
 sky130_fd_sc_hd__a22o_1 _28758_ (.A1(instr_lb),
    .A2(_07774_),
    .B1(_07760_),
    .B2(_07776_),
    .X(_01220_));
 sky130_fd_sc_hd__clkbuf_2 _28759_ (.A(_07706_),
    .X(_07777_));
 sky130_fd_sc_hd__a22o_1 _28760_ (.A1(instr_lh),
    .A2(_07777_),
    .B1(_07764_),
    .B2(_07776_),
    .X(_01221_));
 sky130_fd_sc_hd__nor3b_4 _28761_ (.A(\mem_rdata_q[14] ),
    .B(\mem_rdata_q[12] ),
    .C_N(\mem_rdata_q[13] ),
    .Y(_07778_));
 sky130_fd_sc_hd__a22o_1 _28762_ (.A1(instr_lw),
    .A2(_07777_),
    .B1(_07776_),
    .B2(_07778_),
    .X(_01222_));
 sky130_fd_sc_hd__a22o_1 _28763_ (.A1(instr_lbu),
    .A2(_07777_),
    .B1(_07765_),
    .B2(_07776_),
    .X(_01223_));
 sky130_fd_sc_hd__a22o_1 _28764_ (.A1(instr_lhu),
    .A2(_07777_),
    .B1(_07767_),
    .B2(_07776_),
    .X(_01224_));
 sky130_vsdinv _28765_ (.A(_08519_),
    .Y(_07779_));
 sky130_fd_sc_hd__nand2_1 _28766_ (.A(_07693_),
    .B(_07760_),
    .Y(_07780_));
 sky130_fd_sc_hd__a2bb2o_1 _28767_ (.A1_N(_07779_),
    .A2_N(_07780_),
    .B1(_07774_),
    .B2(instr_sb),
    .X(_01225_));
 sky130_fd_sc_hd__and3_1 _28768_ (.A(_08519_),
    .B(_07739_),
    .C(_07764_),
    .X(_07781_));
 sky130_fd_sc_hd__a21o_1 _28769_ (.A1(instr_sh),
    .A2(_07774_),
    .B1(_07781_),
    .X(_01226_));
 sky130_fd_sc_hd__clkbuf_2 _28770_ (.A(is_alu_reg_imm),
    .X(_07782_));
 sky130_fd_sc_hd__and3_1 _28771_ (.A(_08321_),
    .B(_07782_),
    .C(_07694_),
    .X(_07783_));
 sky130_fd_sc_hd__clkbuf_2 _28772_ (.A(_07783_),
    .X(_07784_));
 sky130_fd_sc_hd__a22o_1 _28773_ (.A1(net453),
    .A2(_07769_),
    .B1(net372),
    .B2(_07784_),
    .X(_01227_));
 sky130_fd_sc_hd__a22o_1 _28774_ (.A1(net472),
    .A2(_07769_),
    .B1(_07778_),
    .B2(_07784_),
    .X(_01228_));
 sky130_fd_sc_hd__and3b_1 _28775_ (.A_N(_07717_),
    .B(_07715_),
    .C(_07713_),
    .X(_07785_));
 sky130_fd_sc_hd__a22o_1 _28776_ (.A1(instr_sltiu),
    .A2(_07769_),
    .B1(_07784_),
    .B2(_07785_),
    .X(_01229_));
 sky130_fd_sc_hd__a22o_1 _28777_ (.A1(net464),
    .A2(_07769_),
    .B1(_07765_),
    .B2(_07784_),
    .X(_01230_));
 sky130_fd_sc_hd__a22o_1 _28778_ (.A1(instr_ori),
    .A2(_07769_),
    .B1(_07768_),
    .B2(_07784_),
    .X(_01231_));
 sky130_fd_sc_hd__clkbuf_2 _28779_ (.A(_07757_),
    .X(_07786_));
 sky130_fd_sc_hd__a22o_1 _28780_ (.A1(net471),
    .A2(_07786_),
    .B1(_07770_),
    .B2(_07784_),
    .X(_01232_));
 sky130_fd_sc_hd__and3_1 _28781_ (.A(_08519_),
    .B(_07695_),
    .C(_07778_),
    .X(_07787_));
 sky130_fd_sc_hd__a21o_1 _28782_ (.A1(instr_sw),
    .A2(_07774_),
    .B1(_07787_),
    .X(_01233_));
 sky130_fd_sc_hd__and2_1 _28783_ (.A(_07782_),
    .B(_07701_),
    .X(_07788_));
 sky130_fd_sc_hd__or4_1 _28784_ (.A(\mem_rdata_q[26] ),
    .B(\mem_rdata_q[27] ),
    .C(\mem_rdata_q[28] ),
    .D(\mem_rdata_q[25] ),
    .X(_07789_));
 sky130_fd_sc_hd__or2_1 _28785_ (.A(\mem_rdata_q[31] ),
    .B(_07742_),
    .X(_07790_));
 sky130_fd_sc_hd__nor2_1 _28786_ (.A(_07745_),
    .B(_07790_),
    .Y(_07791_));
 sky130_fd_sc_hd__and2b_1 _28787_ (.A_N(_07789_),
    .B(_07791_),
    .X(_07792_));
 sky130_fd_sc_hd__and3_1 _28788_ (.A(_07764_),
    .B(_07788_),
    .C(_07792_),
    .X(_07793_));
 sky130_fd_sc_hd__a21o_1 _28789_ (.A1(instr_slli),
    .A2(_07774_),
    .B1(_07793_),
    .X(_01234_));
 sky130_fd_sc_hd__or3_1 _28790_ (.A(\mem_rdata_q[30] ),
    .B(_07789_),
    .C(_07790_),
    .X(_07794_));
 sky130_fd_sc_hd__nor2_2 _28791_ (.A(_07705_),
    .B(_07794_),
    .Y(_07795_));
 sky130_fd_sc_hd__buf_2 _28792_ (.A(_07706_),
    .X(_07796_));
 sky130_fd_sc_hd__a32o_1 _28793_ (.A1(_07782_),
    .A2(_07767_),
    .A3(_07795_),
    .B1(_07796_),
    .B2(net456),
    .X(_01235_));
 sky130_fd_sc_hd__and3_1 _28794_ (.A(_08322_),
    .B(is_alu_reg_reg),
    .C(net372),
    .X(_07797_));
 sky130_fd_sc_hd__a22o_1 _28795_ (.A1(net457),
    .A2(_07786_),
    .B1(_07795_),
    .B2(_07797_),
    .X(_01236_));
 sky130_vsdinv _28796_ (.A(_07745_),
    .Y(_07798_));
 sky130_fd_sc_hd__nor4_1 _28797_ (.A(_07798_),
    .B(_07728_),
    .C(_07789_),
    .D(_07790_),
    .Y(_07799_));
 sky130_fd_sc_hd__a22o_1 _28798_ (.A1(_10430_),
    .A2(_07786_),
    .B1(_07797_),
    .B2(net370),
    .X(_01237_));
 sky130_fd_sc_hd__and3_1 _28799_ (.A(_08321_),
    .B(is_alu_reg_reg),
    .C(_07795_),
    .X(_07800_));
 sky130_fd_sc_hd__clkbuf_2 _28800_ (.A(_07800_),
    .X(_07801_));
 sky130_fd_sc_hd__a22o_1 _28801_ (.A1(instr_sll),
    .A2(_07786_),
    .B1(_07764_),
    .B2(_07801_),
    .X(_01238_));
 sky130_fd_sc_hd__a22o_1 _28802_ (.A1(instr_slt),
    .A2(_07786_),
    .B1(_07778_),
    .B2(_07801_),
    .X(_01239_));
 sky130_fd_sc_hd__a22o_1 _28803_ (.A1(net473),
    .A2(_07786_),
    .B1(_07785_),
    .B2(_07801_),
    .X(_01240_));
 sky130_fd_sc_hd__a22o_1 _28804_ (.A1(instr_xor),
    .A2(_07758_),
    .B1(_07765_),
    .B2(_07801_),
    .X(_01241_));
 sky130_fd_sc_hd__and3_1 _28805_ (.A(_08322_),
    .B(is_alu_reg_reg),
    .C(_07767_),
    .X(_07802_));
 sky130_fd_sc_hd__a22o_1 _28806_ (.A1(net467),
    .A2(_07758_),
    .B1(_07795_),
    .B2(_07802_),
    .X(_01242_));
 sky130_fd_sc_hd__a22o_1 _28807_ (.A1(instr_sra),
    .A2(_07758_),
    .B1(net370),
    .B2(_07802_),
    .X(_01243_));
 sky130_fd_sc_hd__a22o_1 _28808_ (.A1(instr_or),
    .A2(_07758_),
    .B1(_07768_),
    .B2(_07801_),
    .X(_01244_));
 sky130_fd_sc_hd__a22o_1 _28809_ (.A1(net470),
    .A2(_07758_),
    .B1(_07770_),
    .B2(_07801_),
    .X(_01245_));
 sky130_fd_sc_hd__buf_2 _28810_ (.A(_07728_),
    .X(_07803_));
 sky130_fd_sc_hd__a32o_1 _28811_ (.A1(_07782_),
    .A2(_07767_),
    .A3(net370),
    .B1(_07803_),
    .B2(instr_srai),
    .X(_01246_));
 sky130_fd_sc_hd__nor2_1 _28812_ (.A(_07742_),
    .B(\mem_rdata_q[28] ),
    .Y(_07804_));
 sky130_fd_sc_hd__and4_1 _28813_ (.A(_07747_),
    .B(_07745_),
    .C(_07701_),
    .D(_07804_),
    .X(_07805_));
 sky130_fd_sc_hd__nor2_1 _28814_ (.A(_07732_),
    .B(\mem_rdata_q[24] ),
    .Y(_07806_));
 sky130_fd_sc_hd__and4bb_1 _28815_ (.A_N(_07734_),
    .B_N(_07736_),
    .C(_07805_),
    .D(_07806_),
    .X(_07807_));
 sky130_fd_sc_hd__or3_1 _28816_ (.A(\mem_rdata_q[23] ),
    .B(\mem_rdata_q[22] ),
    .C(\mem_rdata_q[21] ),
    .X(_07808_));
 sky130_fd_sc_hd__nand4b_1 _28817_ (.A_N(\mem_rdata_q[3] ),
    .B(\mem_rdata_q[4] ),
    .C(\mem_rdata_q[5] ),
    .D(\mem_rdata_q[6] ),
    .Y(_07809_));
 sky130_fd_sc_hd__or4_1 _28818_ (.A(\mem_rdata_q[17] ),
    .B(\mem_rdata_q[16] ),
    .C(\mem_rdata_q[15] ),
    .D(\mem_rdata_q[2] ),
    .X(_07810_));
 sky130_fd_sc_hd__nand2_1 _28819_ (.A(\mem_rdata_q[0] ),
    .B(\mem_rdata_q[1] ),
    .Y(_07811_));
 sky130_fd_sc_hd__or3_1 _28820_ (.A(\mem_rdata_q[19] ),
    .B(\mem_rdata_q[18] ),
    .C(_07811_),
    .X(_07812_));
 sky130_fd_sc_hd__nor3_1 _28821_ (.A(_07809_),
    .B(_07810_),
    .C(_07812_),
    .Y(_07813_));
 sky130_fd_sc_hd__nand2_1 _28822_ (.A(_07778_),
    .B(_07813_),
    .Y(_07814_));
 sky130_fd_sc_hd__nor2_1 _28823_ (.A(_07808_),
    .B(_07814_),
    .Y(_07815_));
 sky130_fd_sc_hd__a22o_1 _28824_ (.A1(net469),
    .A2(_07777_),
    .B1(_07807_),
    .B2(_07815_),
    .X(_01247_));
 sky130_fd_sc_hd__and4b_1 _28825_ (.A_N(_07734_),
    .B(\mem_rdata_q[27] ),
    .C(_07805_),
    .D(_07806_),
    .X(_07816_));
 sky130_fd_sc_hd__a22o_1 _28826_ (.A1(_08652_),
    .A2(_07777_),
    .B1(_07815_),
    .B2(_07816_),
    .X(_01248_));
 sky130_fd_sc_hd__or4b_1 _28827_ (.A(\mem_rdata_q[23] ),
    .B(\mem_rdata_q[22] ),
    .C(\mem_rdata_q[20] ),
    .D_N(\mem_rdata_q[21] ),
    .X(_07817_));
 sky130_fd_sc_hd__nor2_1 _28828_ (.A(_07814_),
    .B(_07817_),
    .Y(_07818_));
 sky130_fd_sc_hd__a22o_1 _28829_ (.A1(_08749_),
    .A2(_07796_),
    .B1(_07807_),
    .B2(_07818_),
    .X(_01249_));
 sky130_fd_sc_hd__a22o_1 _28830_ (.A1(_08802_),
    .A2(_07796_),
    .B1(_07816_),
    .B2(_07818_),
    .X(_01250_));
 sky130_fd_sc_hd__or3_1 _28831_ (.A(_07809_),
    .B(_07810_),
    .C(_07812_),
    .X(_07819_));
 sky130_fd_sc_hd__or3_1 _28832_ (.A(\mem_rdata_q[7] ),
    .B(\mem_rdata_q[11] ),
    .C(\mem_rdata_q[8] ),
    .X(_07820_));
 sky130_fd_sc_hd__or4_1 _28833_ (.A(\mem_rdata_q[24] ),
    .B(_07780_),
    .C(_07794_),
    .D(_07808_),
    .X(_07821_));
 sky130_fd_sc_hd__or4_1 _28834_ (.A(\mem_rdata_q[10] ),
    .B(\mem_rdata_q[9] ),
    .C(_07820_),
    .D(_07821_),
    .X(_07822_));
 sky130_fd_sc_hd__a2bb2o_1 _28835_ (.A1_N(_07819_),
    .A2_N(_07822_),
    .B1(instr_ecall_ebreak),
    .B2(_07774_),
    .X(_01251_));
 sky130_fd_sc_hd__or3b_1 _28836_ (.A(_07811_),
    .B(\mem_rdata_q[2] ),
    .C_N(\mem_rdata_q[3] ),
    .X(_07823_));
 sky130_fd_sc_hd__nor4_2 _28837_ (.A(\mem_rdata_q[4] ),
    .B(\mem_rdata_q[5] ),
    .C(\mem_rdata_q[6] ),
    .D(_07823_),
    .Y(_07824_));
 sky130_fd_sc_hd__a22o_1 _28838_ (.A1(instr_getq),
    .A2(_07796_),
    .B1(_07795_),
    .B2(_07824_),
    .X(_01252_));
 sky130_fd_sc_hd__and2b_1 _28839_ (.A_N(_07736_),
    .B(_07824_),
    .X(_07825_));
 sky130_fd_sc_hd__and4b_1 _28840_ (.A_N(_07734_),
    .B(_07732_),
    .C(_07741_),
    .D(_07791_),
    .X(_07826_));
 sky130_fd_sc_hd__a22o_1 _28841_ (.A1(instr_setq),
    .A2(_07796_),
    .B1(_07825_),
    .B2(_07826_),
    .X(_01253_));
 sky130_vsdinv _28842_ (.A(_00639_),
    .Y(_07827_));
 sky130_fd_sc_hd__or3_1 _28843_ (.A(_00617_),
    .B(_00618_),
    .C(_00619_),
    .X(_07828_));
 sky130_fd_sc_hd__nand3b_1 _28844_ (.A_N(_00615_),
    .B(_00614_),
    .C(_00613_),
    .Y(_07829_));
 sky130_fd_sc_hd__or4b_1 _28845_ (.A(_00638_),
    .B(_00642_),
    .C(_00643_),
    .D_N(_00616_),
    .X(_07830_));
 sky130_fd_sc_hd__or4_1 _28846_ (.A(_00644_),
    .B(_07828_),
    .C(_07829_),
    .D(_07830_),
    .X(_07831_));
 sky130_fd_sc_hd__or3_1 _28847_ (.A(_00640_),
    .B(_00641_),
    .C(_07831_),
    .X(_07832_));
 sky130_fd_sc_hd__nor2_2 _28848_ (.A(_07827_),
    .B(_07832_),
    .Y(_07833_));
 sky130_fd_sc_hd__clkbuf_4 _28849_ (.A(_05512_),
    .X(_07834_));
 sky130_fd_sc_hd__mux2_1 _28850_ (.A0(instr_retirq),
    .A1(_07833_),
    .S(_07834_),
    .X(_07835_));
 sky130_fd_sc_hd__clkbuf_1 _28851_ (.A(_07835_),
    .X(_01254_));
 sky130_fd_sc_hd__and4_1 _28852_ (.A(_07734_),
    .B(_07732_),
    .C(_07741_),
    .D(_07791_),
    .X(_07836_));
 sky130_fd_sc_hd__a22o_1 _28853_ (.A1(_08639_),
    .A2(_07796_),
    .B1(_07825_),
    .B2(_07836_),
    .X(_01255_));
 sky130_fd_sc_hd__nor4_1 _28854_ (.A(_08536_),
    .B(_00639_),
    .C(_00641_),
    .D(_07831_),
    .Y(_07837_));
 sky130_fd_sc_hd__a22o_1 _28855_ (.A1(_08207_),
    .A2(_07771_),
    .B1(_00640_),
    .B2(_07837_),
    .X(_01256_));
 sky130_fd_sc_hd__and2_1 _28856_ (.A(_08643_),
    .B(_07706_),
    .X(_07838_));
 sky130_fd_sc_hd__a31o_1 _28857_ (.A1(_07736_),
    .A2(_07824_),
    .A3(_07826_),
    .B1(_07838_),
    .X(_01257_));
 sky130_fd_sc_hd__a2bb2o_1 _28858_ (.A1_N(_07833_),
    .A2_N(_05540_),
    .B1(_05536_),
    .B2(\decoded_rs1[0] ),
    .X(_01258_));
 sky130_fd_sc_hd__a2bb2o_1 _28859_ (.A1_N(_07833_),
    .A2_N(_05542_),
    .B1(_05536_),
    .B2(\decoded_rs1[1] ),
    .X(_01259_));
 sky130_fd_sc_hd__a2bb2o_1 _28860_ (.A1_N(_07833_),
    .A2_N(_05544_),
    .B1(_07749_),
    .B2(\decoded_rs1[2] ),
    .X(_01260_));
 sky130_fd_sc_hd__a2bb2o_1 _28861_ (.A1_N(_07833_),
    .A2_N(_05546_),
    .B1(_07749_),
    .B2(\decoded_rs1[3] ),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _28862_ (.A0(\decoded_rd[0] ),
    .A1(_00620_),
    .S(_07834_),
    .X(_07839_));
 sky130_fd_sc_hd__clkbuf_1 _28863_ (.A(_07839_),
    .X(_01262_));
 sky130_fd_sc_hd__mux2_1 _28864_ (.A0(\decoded_rd[1] ),
    .A1(_00621_),
    .S(_07834_),
    .X(_07840_));
 sky130_fd_sc_hd__clkbuf_1 _28865_ (.A(_07840_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _28866_ (.A0(\decoded_rd[2] ),
    .A1(_00622_),
    .S(_07834_),
    .X(_07841_));
 sky130_fd_sc_hd__clkbuf_1 _28867_ (.A(_07841_),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _28868_ (.A0(\decoded_rd[3] ),
    .A1(_00623_),
    .S(_07834_),
    .X(_07842_));
 sky130_fd_sc_hd__clkbuf_1 _28869_ (.A(_07842_),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _28870_ (.A0(\decoded_rd[4] ),
    .A1(_00624_),
    .S(_07834_),
    .X(_07843_));
 sky130_fd_sc_hd__clkbuf_1 _28871_ (.A(_07843_),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _28872_ (.A0(_08554_),
    .A1(_00633_),
    .S(_05537_),
    .X(_07844_));
 sky130_fd_sc_hd__clkbuf_1 _28873_ (.A(_07844_),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_2 _28874_ (.A0(_08546_),
    .A1(_00634_),
    .S(_05537_),
    .X(_07845_));
 sky130_fd_sc_hd__clkbuf_1 _28875_ (.A(_07845_),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _28876_ (.A0(\decoded_imm_uj[2] ),
    .A1(_00635_),
    .S(_05537_),
    .X(_07846_));
 sky130_fd_sc_hd__clkbuf_1 _28877_ (.A(_07846_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _28878_ (.A0(\decoded_imm_uj[3] ),
    .A1(_00636_),
    .S(_05537_),
    .X(_07847_));
 sky130_fd_sc_hd__clkbuf_1 _28879_ (.A(_07847_),
    .X(_01270_));
 sky130_fd_sc_hd__and3_1 _28880_ (.A(is_sb_sh_sw),
    .B(\mem_rdata_q[7] ),
    .C(_07743_),
    .X(_07848_));
 sky130_fd_sc_hd__or3_2 _28881_ (.A(instr_jalr),
    .B(is_lb_lh_lw_lbu_lhu),
    .C(is_alu_reg_imm),
    .X(_07849_));
 sky130_fd_sc_hd__buf_1 _28882_ (.A(_07849_),
    .X(_07850_));
 sky130_fd_sc_hd__and3_1 _28883_ (.A(\mem_rdata_q[20] ),
    .B(_07743_),
    .C(_07850_),
    .X(_07851_));
 sky130_fd_sc_hd__a211o_1 _28884_ (.A1(_08668_),
    .A2(_07803_),
    .B1(_07848_),
    .C1(_07851_),
    .X(_01271_));
 sky130_fd_sc_hd__nor2_1 _28885_ (.A(_00616_),
    .B(_07829_),
    .Y(_07852_));
 sky130_fd_sc_hd__nor2_1 _28886_ (.A(_08536_),
    .B(_07828_),
    .Y(_07853_));
 sky130_fd_sc_hd__a22o_1 _28887_ (.A1(is_lb_lh_lw_lbu_lhu),
    .A2(_07771_),
    .B1(_07852_),
    .B2(_07853_),
    .X(_01272_));
 sky130_fd_sc_hd__or4b_1 _28888_ (.A(_07747_),
    .B(_07789_),
    .C(_07742_),
    .D_N(_07767_),
    .X(_07854_));
 sky130_vsdinv _28889_ (.A(_07854_),
    .Y(_07855_));
 sky130_fd_sc_hd__a221o_1 _28890_ (.A1(_07385_),
    .A2(_07803_),
    .B1(_07788_),
    .B2(_07855_),
    .C1(_07793_),
    .X(_01273_));
 sky130_fd_sc_hd__a211o_1 _28891_ (.A1(_07782_),
    .A2(_07763_),
    .B1(_07706_),
    .C1(instr_jalr),
    .X(_07856_));
 sky130_fd_sc_hd__o21a_1 _28892_ (.A1(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .A2(_07740_),
    .B1(_07856_),
    .X(_01274_));
 sky130_fd_sc_hd__and3b_1 _28893_ (.A_N(_00617_),
    .B(_00618_),
    .C(_07852_),
    .X(_07857_));
 sky130_fd_sc_hd__a22o_1 _28894_ (.A1(_08519_),
    .A2(_07771_),
    .B1(_07752_),
    .B2(_07857_),
    .X(_01275_));
 sky130_fd_sc_hd__and3_1 _28895_ (.A(_05513_),
    .B(_00619_),
    .C(_07857_),
    .X(_07858_));
 sky130_fd_sc_hd__a31o_1 _28896_ (.A1(_08294_),
    .A2(_06184_),
    .A3(_07749_),
    .B1(_07858_),
    .X(_01276_));
 sky130_fd_sc_hd__a22o_1 _28897_ (.A1(_07782_),
    .A2(_07771_),
    .B1(_07754_),
    .B2(_07852_),
    .X(_01277_));
 sky130_fd_sc_hd__a22o_1 _28898_ (.A1(is_alu_reg_reg),
    .A2(_07771_),
    .B1(_07753_),
    .B2(_07852_),
    .X(_01278_));
 sky130_fd_sc_hd__o21a_1 _28899_ (.A1(_08294_),
    .A2(_08219_),
    .B1(_07759_),
    .X(_01279_));
 sky130_fd_sc_hd__nand2_1 _28900_ (.A(_10320_),
    .B(_05748_),
    .Y(_07859_));
 sky130_fd_sc_hd__clkbuf_4 _28901_ (.A(_05745_),
    .X(_07860_));
 sky130_fd_sc_hd__o21ba_2 _28902_ (.A1(_08525_),
    .A2(_05738_),
    .B1_N(_07860_),
    .X(_07861_));
 sky130_fd_sc_hd__a2bb2o_1 _28903_ (.A1_N(_08163_),
    .A2_N(_07859_),
    .B1(_07861_),
    .B2(net129),
    .X(_01280_));
 sky130_fd_sc_hd__nand2_1 _28904_ (.A(\mem_state[0] ),
    .B(_05737_),
    .Y(_07862_));
 sky130_fd_sc_hd__or4_1 _28905_ (.A(_08151_),
    .B(_08522_),
    .C(\mem_state[1] ),
    .D(_07862_),
    .X(_07863_));
 sky130_fd_sc_hd__o21ai_1 _28906_ (.A1(_05738_),
    .A2(_05739_),
    .B1(_07863_),
    .Y(_07864_));
 sky130_fd_sc_hd__or3b_1 _28907_ (.A(_05738_),
    .B(_08522_),
    .C_N(_08156_),
    .X(_07865_));
 sky130_fd_sc_hd__o211a_1 _28908_ (.A1(_05738_),
    .A2(_05741_),
    .B1(_05742_),
    .C1(_07865_),
    .X(_07866_));
 sky130_fd_sc_hd__mux2_1 _28909_ (.A0(\mem_state[0] ),
    .A1(_07864_),
    .S(_07866_),
    .X(_07867_));
 sky130_fd_sc_hd__clkbuf_1 _28910_ (.A(_07867_),
    .X(_01281_));
 sky130_fd_sc_hd__or2b_1 _28911_ (.A(_07860_),
    .B_N(_07863_),
    .X(_07868_));
 sky130_fd_sc_hd__mux2_1 _28912_ (.A0(\mem_state[1] ),
    .A1(_07868_),
    .S(_07866_),
    .X(_07869_));
 sky130_fd_sc_hd__clkbuf_1 _28913_ (.A(_07869_),
    .X(_01282_));
 sky130_fd_sc_hd__clkbuf_2 _28914_ (.A(_07860_),
    .X(_07870_));
 sky130_fd_sc_hd__mux2_1 _28915_ (.A0(net199),
    .A1(_10270_),
    .S(_07870_),
    .X(_07871_));
 sky130_fd_sc_hd__clkbuf_1 _28916_ (.A(_07871_),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _28917_ (.A0(net210),
    .A1(_10108_),
    .S(_07870_),
    .X(_07872_));
 sky130_fd_sc_hd__clkbuf_1 _28918_ (.A(_07872_),
    .X(_01284_));
 sky130_fd_sc_hd__clkbuf_2 _28919_ (.A(_07860_),
    .X(_07873_));
 sky130_fd_sc_hd__mux2_1 _28920_ (.A0(net221),
    .A1(_10273_),
    .S(_07873_),
    .X(_07874_));
 sky130_fd_sc_hd__clkbuf_1 _28921_ (.A(_07874_),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _28922_ (.A0(net224),
    .A1(_04961_),
    .S(_07873_),
    .X(_07875_));
 sky130_fd_sc_hd__clkbuf_1 _28923_ (.A(_07875_),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _28924_ (.A0(net225),
    .A1(_04755_),
    .S(_07873_),
    .X(_07876_));
 sky130_fd_sc_hd__clkbuf_1 _28925_ (.A(_07876_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _28926_ (.A0(net226),
    .A1(_10277_),
    .S(_07873_),
    .X(_07877_));
 sky130_fd_sc_hd__clkbuf_1 _28927_ (.A(_07877_),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _28928_ (.A0(net227),
    .A1(_10279_),
    .S(_07873_),
    .X(_07878_));
 sky130_fd_sc_hd__clkbuf_1 _28929_ (.A(_07878_),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _28930_ (.A0(net228),
    .A1(_10280_),
    .S(_07873_),
    .X(_07879_));
 sky130_fd_sc_hd__clkbuf_1 _28931_ (.A(_07879_),
    .X(_01290_));
 sky130_fd_sc_hd__clkbuf_2 _28932_ (.A(_07860_),
    .X(_07880_));
 sky130_fd_sc_hd__mux2_1 _28933_ (.A0(net229),
    .A1(net191),
    .S(_07880_),
    .X(_07881_));
 sky130_fd_sc_hd__clkbuf_1 _28934_ (.A(_07881_),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _28935_ (.A0(net230),
    .A1(net192),
    .S(_07880_),
    .X(_07882_));
 sky130_fd_sc_hd__clkbuf_1 _28936_ (.A(_07882_),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _28937_ (.A0(net200),
    .A1(net162),
    .S(_07880_),
    .X(_07883_));
 sky130_fd_sc_hd__clkbuf_1 _28938_ (.A(_07883_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _28939_ (.A0(net201),
    .A1(net163),
    .S(_07880_),
    .X(_07884_));
 sky130_fd_sc_hd__clkbuf_1 _28940_ (.A(_07884_),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _28941_ (.A0(net202),
    .A1(net164),
    .S(_07880_),
    .X(_07885_));
 sky130_fd_sc_hd__clkbuf_1 _28942_ (.A(_07885_),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _28943_ (.A0(net203),
    .A1(net165),
    .S(_07880_),
    .X(_07886_));
 sky130_fd_sc_hd__clkbuf_1 _28944_ (.A(_07886_),
    .X(_01296_));
 sky130_fd_sc_hd__buf_2 _28945_ (.A(_07860_),
    .X(_07887_));
 sky130_fd_sc_hd__mux2_1 _28946_ (.A0(net204),
    .A1(net166),
    .S(_07887_),
    .X(_07888_));
 sky130_fd_sc_hd__clkbuf_1 _28947_ (.A(_07888_),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _28948_ (.A0(net205),
    .A1(net167),
    .S(_07887_),
    .X(_07889_));
 sky130_fd_sc_hd__clkbuf_1 _28949_ (.A(_07889_),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _28950_ (.A0(net206),
    .A1(net168),
    .S(_07887_),
    .X(_07890_));
 sky130_fd_sc_hd__clkbuf_1 _28951_ (.A(_07890_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _28952_ (.A0(net207),
    .A1(net169),
    .S(_07887_),
    .X(_07891_));
 sky130_fd_sc_hd__clkbuf_1 _28953_ (.A(_07891_),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _28954_ (.A0(net208),
    .A1(net170),
    .S(_07887_),
    .X(_07892_));
 sky130_fd_sc_hd__clkbuf_1 _28955_ (.A(_07892_),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _28956_ (.A0(net209),
    .A1(net171),
    .S(_07887_),
    .X(_07893_));
 sky130_fd_sc_hd__clkbuf_1 _28957_ (.A(_07893_),
    .X(_01302_));
 sky130_fd_sc_hd__clkbuf_4 _28958_ (.A(_05745_),
    .X(_07894_));
 sky130_fd_sc_hd__mux2_1 _28959_ (.A0(net211),
    .A1(net173),
    .S(_07894_),
    .X(_07895_));
 sky130_fd_sc_hd__clkbuf_1 _28960_ (.A(_07895_),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _28961_ (.A0(net212),
    .A1(net174),
    .S(_07894_),
    .X(_07896_));
 sky130_fd_sc_hd__clkbuf_1 _28962_ (.A(_07896_),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _28963_ (.A0(net213),
    .A1(net175),
    .S(_07894_),
    .X(_07897_));
 sky130_fd_sc_hd__clkbuf_1 _28964_ (.A(_07897_),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _28965_ (.A0(net214),
    .A1(net176),
    .S(_07894_),
    .X(_07898_));
 sky130_fd_sc_hd__clkbuf_1 _28966_ (.A(_07898_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _28967_ (.A0(net215),
    .A1(net177),
    .S(_07894_),
    .X(_07899_));
 sky130_fd_sc_hd__clkbuf_1 _28968_ (.A(_07899_),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _28969_ (.A0(net216),
    .A1(net178),
    .S(_07894_),
    .X(_07900_));
 sky130_fd_sc_hd__clkbuf_1 _28970_ (.A(_07900_),
    .X(_01308_));
 sky130_fd_sc_hd__buf_2 _28971_ (.A(_05745_),
    .X(_07901_));
 sky130_fd_sc_hd__mux2_1 _28972_ (.A0(net217),
    .A1(net179),
    .S(_07901_),
    .X(_07902_));
 sky130_fd_sc_hd__clkbuf_1 _28973_ (.A(_07902_),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _28974_ (.A0(net218),
    .A1(net180),
    .S(_07901_),
    .X(_07903_));
 sky130_fd_sc_hd__clkbuf_1 _28975_ (.A(_07903_),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _28976_ (.A0(net219),
    .A1(net181),
    .S(_07901_),
    .X(_07904_));
 sky130_fd_sc_hd__clkbuf_1 _28977_ (.A(_07904_),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _28978_ (.A0(net220),
    .A1(net182),
    .S(_07901_),
    .X(_07905_));
 sky130_fd_sc_hd__clkbuf_1 _28979_ (.A(_07905_),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _28980_ (.A0(net222),
    .A1(net184),
    .S(_07901_),
    .X(_07906_));
 sky130_fd_sc_hd__clkbuf_1 _28981_ (.A(_07906_),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _28982_ (.A0(net223),
    .A1(net185),
    .S(_07901_),
    .X(_07907_));
 sky130_fd_sc_hd__clkbuf_1 _28983_ (.A(_07907_),
    .X(_01314_));
 sky130_fd_sc_hd__a32o_1 _28984_ (.A1(_08525_),
    .A2(net194),
    .A3(_07870_),
    .B1(_07861_),
    .B2(net231),
    .X(_01315_));
 sky130_fd_sc_hd__a32o_1 _28985_ (.A1(_08525_),
    .A2(net195),
    .A3(_07870_),
    .B1(_07861_),
    .B2(net232),
    .X(_01316_));
 sky130_fd_sc_hd__a32o_1 _28986_ (.A1(_08525_),
    .A2(net196),
    .A3(_07870_),
    .B1(_07861_),
    .B2(net233),
    .X(_01317_));
 sky130_fd_sc_hd__a32o_1 _28987_ (.A1(_08525_),
    .A2(net197),
    .A3(_07870_),
    .B1(_07861_),
    .B2(net234),
    .X(_01318_));
 sky130_fd_sc_hd__and2b_1 _28988_ (.A_N(_04773_),
    .B(_04709_),
    .X(_07908_));
 sky130_fd_sc_hd__clkbuf_1 _28989_ (.A(_07908_),
    .X(_01319_));
 sky130_fd_sc_hd__and2b_1 _28990_ (.A_N(_04773_),
    .B(_04727_),
    .X(_07909_));
 sky130_fd_sc_hd__clkbuf_1 _28991_ (.A(_07909_),
    .X(_01320_));
 sky130_fd_sc_hd__and2b_1 _28992_ (.A_N(_04773_),
    .B(_04740_),
    .X(_07910_));
 sky130_fd_sc_hd__clkbuf_1 _28993_ (.A(_07910_),
    .X(_01321_));
 sky130_fd_sc_hd__and2b_1 _28994_ (.A_N(_04773_),
    .B(_04752_),
    .X(_07911_));
 sky130_fd_sc_hd__clkbuf_1 _28995_ (.A(_07911_),
    .X(_01322_));
 sky130_fd_sc_hd__clkbuf_2 _28996_ (.A(_04815_),
    .X(_07912_));
 sky130_fd_sc_hd__nor3_1 _28997_ (.A(_07397_),
    .B(_07912_),
    .C(_04760_),
    .Y(_01323_));
 sky130_fd_sc_hd__and2b_1 _28998_ (.A_N(_04773_),
    .B(_04781_),
    .X(_07913_));
 sky130_fd_sc_hd__clkbuf_1 _28999_ (.A(_07913_),
    .X(_01324_));
 sky130_fd_sc_hd__and2b_1 _29000_ (.A_N(_04946_),
    .B(_04791_),
    .X(_07914_));
 sky130_fd_sc_hd__clkbuf_1 _29001_ (.A(_07914_),
    .X(_01325_));
 sky130_fd_sc_hd__and2b_1 _29002_ (.A_N(_04946_),
    .B(_04798_),
    .X(_07915_));
 sky130_fd_sc_hd__clkbuf_1 _29003_ (.A(_07915_),
    .X(_01326_));
 sky130_fd_sc_hd__nor2_1 _29004_ (.A(_04763_),
    .B(_04695_),
    .Y(_07916_));
 sky130_fd_sc_hd__a211oi_1 _29005_ (.A1(_07397_),
    .A2(_04708_),
    .B1(_07916_),
    .C1(_07912_),
    .Y(_01327_));
 sky130_fd_sc_hd__nor2_1 _29006_ (.A(_04763_),
    .B(_04715_),
    .Y(_07917_));
 sky130_fd_sc_hd__a211oi_1 _29007_ (.A1(_07397_),
    .A2(_04726_),
    .B1(_07917_),
    .C1(_07912_),
    .Y(_01328_));
 sky130_fd_sc_hd__nor2_1 _29008_ (.A(_04763_),
    .B(_04735_),
    .Y(_07918_));
 sky130_fd_sc_hd__a211oi_1 _29009_ (.A1(_07397_),
    .A2(_04739_),
    .B1(_07918_),
    .C1(_07912_),
    .Y(_01329_));
 sky130_fd_sc_hd__nor2_1 _29010_ (.A(_04763_),
    .B(_04744_),
    .Y(_07919_));
 sky130_fd_sc_hd__a211oi_1 _29011_ (.A1(_07397_),
    .A2(_04751_),
    .B1(_07919_),
    .C1(_07912_),
    .Y(_01330_));
 sky130_fd_sc_hd__mux2_1 _29012_ (.A0(_04767_),
    .A1(_04760_),
    .S(_04705_),
    .X(_07920_));
 sky130_fd_sc_hd__nor2_1 _29013_ (.A(_04756_),
    .B(_07920_),
    .Y(_01331_));
 sky130_fd_sc_hd__nor2_1 _29014_ (.A(_04961_),
    .B(_04777_),
    .Y(_07921_));
 sky130_fd_sc_hd__a211oi_1 _29015_ (.A1(_04763_),
    .A2(_04780_),
    .B1(_07921_),
    .C1(_07912_),
    .Y(_01332_));
 sky130_fd_sc_hd__and2b_1 _29016_ (.A_N(_04946_),
    .B(_04834_),
    .X(_07922_));
 sky130_fd_sc_hd__clkbuf_1 _29017_ (.A(_07922_),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _29018_ (.A0(_04795_),
    .A1(_04797_),
    .S(_10274_),
    .X(_07923_));
 sky130_fd_sc_hd__and2b_1 _29019_ (.A_N(_04946_),
    .B(_07923_),
    .X(_07924_));
 sky130_fd_sc_hd__clkbuf_1 _29020_ (.A(_07924_),
    .X(_01334_));
 sky130_fd_sc_hd__and2_1 _29021_ (.A(_08216_),
    .B(_07701_),
    .X(_07925_));
 sky130_fd_sc_hd__clkbuf_2 _29022_ (.A(_07925_),
    .X(_07926_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29023_ (.A(_07728_),
    .X(_07927_));
 sky130_fd_sc_hd__and2_1 _29024_ (.A(\decoded_imm[31] ),
    .B(_07927_),
    .X(_07928_));
 sky130_fd_sc_hd__or2_2 _29025_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .B(is_sb_sh_sw),
    .X(_07929_));
 sky130_fd_sc_hd__and2_1 _29026_ (.A(\mem_rdata_q[31] ),
    .B(_07929_),
    .X(_07930_));
 sky130_fd_sc_hd__a22o_1 _29027_ (.A1(_06726_),
    .A2(_05552_),
    .B1(_07849_),
    .B2(\mem_rdata_q[31] ),
    .X(_07931_));
 sky130_fd_sc_hd__o21a_1 _29028_ (.A1(_07930_),
    .A2(_07931_),
    .B1(_07694_),
    .X(_07932_));
 sky130_fd_sc_hd__clkbuf_2 _29029_ (.A(_07932_),
    .X(_07933_));
 sky130_fd_sc_hd__a211o_1 _29030_ (.A1(_07747_),
    .A2(_07926_),
    .B1(_07928_),
    .C1(_07933_),
    .X(_01335_));
 sky130_fd_sc_hd__clkbuf_2 _29031_ (.A(_07925_),
    .X(_07934_));
 sky130_fd_sc_hd__clkbuf_2 _29032_ (.A(_07932_),
    .X(_07935_));
 sky130_fd_sc_hd__a221o_1 _29033_ (.A1(\decoded_imm[30] ),
    .A2(_07803_),
    .B1(_07934_),
    .B2(_07745_),
    .C1(_07935_),
    .X(_01336_));
 sky130_fd_sc_hd__and2_1 _29034_ (.A(\decoded_imm[29] ),
    .B(_07927_),
    .X(_07936_));
 sky130_fd_sc_hd__a211o_1 _29035_ (.A1(_07742_),
    .A2(_07926_),
    .B1(_07936_),
    .C1(_07933_),
    .X(_01337_));
 sky130_fd_sc_hd__and2_1 _29036_ (.A(\decoded_imm[28] ),
    .B(_07927_),
    .X(_07937_));
 sky130_fd_sc_hd__a211o_1 _29037_ (.A1(net454),
    .A2(_07926_),
    .B1(_07937_),
    .C1(_07933_),
    .X(_01338_));
 sky130_fd_sc_hd__and2_1 _29038_ (.A(\decoded_imm[27] ),
    .B(_07927_),
    .X(_07938_));
 sky130_fd_sc_hd__a211o_1 _29039_ (.A1(_07736_),
    .A2(_07926_),
    .B1(_07938_),
    .C1(_07933_),
    .X(_01339_));
 sky130_fd_sc_hd__a221o_1 _29040_ (.A1(\decoded_imm[26] ),
    .A2(_07803_),
    .B1(_07934_),
    .B2(_07734_),
    .C1(_07935_),
    .X(_01340_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29041_ (.A(_07705_),
    .X(_07939_));
 sky130_fd_sc_hd__and2_1 _29042_ (.A(\decoded_imm[25] ),
    .B(_07939_),
    .X(_07940_));
 sky130_fd_sc_hd__a211o_1 _29043_ (.A1(_07732_),
    .A2(_07926_),
    .B1(_07940_),
    .C1(_07933_),
    .X(_01341_));
 sky130_fd_sc_hd__and2_1 _29044_ (.A(\decoded_imm[24] ),
    .B(_07939_),
    .X(_07941_));
 sky130_fd_sc_hd__a211o_1 _29045_ (.A1(\mem_rdata_q[24] ),
    .A2(_07926_),
    .B1(_07941_),
    .C1(_07933_),
    .X(_01342_));
 sky130_fd_sc_hd__and2_1 _29046_ (.A(_09751_),
    .B(_07939_),
    .X(_07942_));
 sky130_fd_sc_hd__a211o_1 _29047_ (.A1(\mem_rdata_q[23] ),
    .A2(_07934_),
    .B1(_07942_),
    .C1(_07935_),
    .X(_01343_));
 sky130_fd_sc_hd__and2_1 _29048_ (.A(\decoded_imm[22] ),
    .B(_07939_),
    .X(_07943_));
 sky130_fd_sc_hd__a211o_1 _29049_ (.A1(\mem_rdata_q[22] ),
    .A2(_07934_),
    .B1(_07943_),
    .C1(_07935_),
    .X(_01344_));
 sky130_fd_sc_hd__and2_1 _29050_ (.A(\decoded_imm[21] ),
    .B(_07939_),
    .X(_07944_));
 sky130_fd_sc_hd__a211o_1 _29051_ (.A1(\mem_rdata_q[21] ),
    .A2(_07934_),
    .B1(_07944_),
    .C1(_07935_),
    .X(_01345_));
 sky130_fd_sc_hd__a221o_1 _29052_ (.A1(\decoded_imm[20] ),
    .A2(_07803_),
    .B1(_07934_),
    .B2(\mem_rdata_q[20] ),
    .C1(_07935_),
    .X(_01346_));
 sky130_fd_sc_hd__a21o_1 _29053_ (.A1(_07747_),
    .A2(_07850_),
    .B1(_07728_),
    .X(_07945_));
 sky130_fd_sc_hd__clkbuf_2 _29054_ (.A(_07945_),
    .X(_07946_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29055_ (.A(_08216_),
    .X(_07947_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29056_ (.A(_07930_),
    .X(_07948_));
 sky130_fd_sc_hd__a221o_1 _29057_ (.A1(_07535_),
    .A2(\decoded_imm_uj[19] ),
    .B1(_07947_),
    .B2(\mem_rdata_q[19] ),
    .C1(_07948_),
    .X(_07949_));
 sky130_fd_sc_hd__o22a_1 _29058_ (.A1(\decoded_imm[19] ),
    .A2(_07740_),
    .B1(_07946_),
    .B2(_07949_),
    .X(_01347_));
 sky130_fd_sc_hd__a221o_1 _29059_ (.A1(_07535_),
    .A2(\decoded_imm_uj[18] ),
    .B1(_07947_),
    .B2(\mem_rdata_q[18] ),
    .C1(_07948_),
    .X(_07950_));
 sky130_fd_sc_hd__o22a_1 _29060_ (.A1(\decoded_imm[18] ),
    .A2(_07740_),
    .B1(_07946_),
    .B2(_07950_),
    .X(_01348_));
 sky130_fd_sc_hd__a221o_1 _29061_ (.A1(_07535_),
    .A2(\decoded_imm_uj[17] ),
    .B1(_07947_),
    .B2(\mem_rdata_q[17] ),
    .C1(_07948_),
    .X(_07951_));
 sky130_fd_sc_hd__o22a_1 _29062_ (.A1(\decoded_imm[17] ),
    .A2(_07740_),
    .B1(_07946_),
    .B2(_07951_),
    .X(_01349_));
 sky130_fd_sc_hd__a221o_1 _29063_ (.A1(_07535_),
    .A2(\decoded_imm_uj[16] ),
    .B1(_07947_),
    .B2(\mem_rdata_q[16] ),
    .C1(_07948_),
    .X(_07952_));
 sky130_fd_sc_hd__o22a_1 _29064_ (.A1(\decoded_imm[16] ),
    .A2(_07740_),
    .B1(_07946_),
    .B2(_07952_),
    .X(_01350_));
 sky130_fd_sc_hd__clkbuf_2 _29065_ (.A(_07739_),
    .X(_07953_));
 sky130_fd_sc_hd__clkbuf_2 _29066_ (.A(_06555_),
    .X(_07954_));
 sky130_fd_sc_hd__a221o_1 _29067_ (.A1(_07954_),
    .A2(\decoded_imm_uj[15] ),
    .B1(_07947_),
    .B2(\mem_rdata_q[15] ),
    .C1(_07948_),
    .X(_07955_));
 sky130_fd_sc_hd__o22a_1 _29068_ (.A1(\decoded_imm[15] ),
    .A2(_07953_),
    .B1(_07946_),
    .B2(_07955_),
    .X(_01351_));
 sky130_fd_sc_hd__a221o_1 _29069_ (.A1(_07954_),
    .A2(\decoded_imm_uj[14] ),
    .B1(_07947_),
    .B2(_07717_),
    .C1(_07948_),
    .X(_07956_));
 sky130_fd_sc_hd__o22a_1 _29070_ (.A1(\decoded_imm[14] ),
    .A2(_07953_),
    .B1(_07946_),
    .B2(_07956_),
    .X(_01352_));
 sky130_fd_sc_hd__a221o_1 _29071_ (.A1(_07954_),
    .A2(\decoded_imm_uj[13] ),
    .B1(_08216_),
    .B2(_07715_),
    .C1(_07930_),
    .X(_07957_));
 sky130_fd_sc_hd__o22a_1 _29072_ (.A1(\decoded_imm[13] ),
    .A2(_07953_),
    .B1(_07945_),
    .B2(_07957_),
    .X(_01353_));
 sky130_fd_sc_hd__a221o_1 _29073_ (.A1(_07954_),
    .A2(\decoded_imm_uj[12] ),
    .B1(_08216_),
    .B2(_07713_),
    .C1(_07930_),
    .X(_07958_));
 sky130_fd_sc_hd__o22a_1 _29074_ (.A1(_09305_),
    .A2(_07953_),
    .B1(_07945_),
    .B2(_07958_),
    .X(_01354_));
 sky130_fd_sc_hd__a22o_1 _29075_ (.A1(_08294_),
    .A2(\mem_rdata_q[7] ),
    .B1(_08554_),
    .B2(_06455_),
    .X(_07959_));
 sky130_fd_sc_hd__a21o_1 _29076_ (.A1(_08519_),
    .A2(_07747_),
    .B1(_07959_),
    .X(_07960_));
 sky130_fd_sc_hd__o22a_1 _29077_ (.A1(\decoded_imm[11] ),
    .A2(_07953_),
    .B1(_07945_),
    .B2(_07960_),
    .X(_01355_));
 sky130_fd_sc_hd__clkbuf_2 _29078_ (.A(_07939_),
    .X(_07961_));
 sky130_fd_sc_hd__nor2_2 _29079_ (.A(decoder_pseudo_trigger),
    .B(_06542_),
    .Y(_07962_));
 sky130_fd_sc_hd__or2_1 _29080_ (.A(_07849_),
    .B(_07929_),
    .X(_07963_));
 sky130_fd_sc_hd__and3_1 _29081_ (.A(_07745_),
    .B(_07743_),
    .C(_07963_),
    .X(_07964_));
 sky130_fd_sc_hd__a221o_1 _29082_ (.A1(_09219_),
    .A2(_07961_),
    .B1(_07962_),
    .B2(\decoded_imm_uj[10] ),
    .C1(_07964_),
    .X(_01356_));
 sky130_fd_sc_hd__and3_1 _29083_ (.A(_07742_),
    .B(_07738_),
    .C(_07963_),
    .X(_07965_));
 sky130_fd_sc_hd__a221o_1 _29084_ (.A1(\decoded_imm[9] ),
    .A2(_07961_),
    .B1(_07962_),
    .B2(\decoded_imm_uj[9] ),
    .C1(_07965_),
    .X(_01357_));
 sky130_fd_sc_hd__and3_1 _29085_ (.A(\mem_rdata_q[28] ),
    .B(_07738_),
    .C(_07963_),
    .X(_07966_));
 sky130_fd_sc_hd__a221o_1 _29086_ (.A1(\decoded_imm[8] ),
    .A2(_07961_),
    .B1(_07962_),
    .B2(\decoded_imm_uj[8] ),
    .C1(_07966_),
    .X(_01358_));
 sky130_fd_sc_hd__and3_1 _29087_ (.A(_07736_),
    .B(_07738_),
    .C(_07963_),
    .X(_07967_));
 sky130_fd_sc_hd__a221o_1 _29088_ (.A1(\decoded_imm[7] ),
    .A2(_07961_),
    .B1(_07962_),
    .B2(\decoded_imm_uj[7] ),
    .C1(_07967_),
    .X(_01359_));
 sky130_fd_sc_hd__and3_1 _29089_ (.A(\mem_rdata_q[26] ),
    .B(_07738_),
    .C(_07963_),
    .X(_07968_));
 sky130_fd_sc_hd__a221o_1 _29090_ (.A1(\decoded_imm[6] ),
    .A2(_07961_),
    .B1(_07962_),
    .B2(\decoded_imm_uj[6] ),
    .C1(_07968_),
    .X(_01360_));
 sky130_fd_sc_hd__and3_1 _29091_ (.A(_07732_),
    .B(_07738_),
    .C(_07963_),
    .X(_07969_));
 sky130_fd_sc_hd__a221o_1 _29092_ (.A1(\decoded_imm[5] ),
    .A2(_07961_),
    .B1(_07962_),
    .B2(\decoded_imm_uj[5] ),
    .C1(_07969_),
    .X(_01361_));
 sky130_fd_sc_hd__and2_1 _29093_ (.A(\mem_rdata_q[24] ),
    .B(_07850_),
    .X(_07970_));
 sky130_fd_sc_hd__a221o_1 _29094_ (.A1(_07954_),
    .A2(\decoded_imm_uj[4] ),
    .B1(_07929_),
    .B2(\mem_rdata_q[11] ),
    .C1(_07729_),
    .X(_07971_));
 sky130_fd_sc_hd__o22a_1 _29095_ (.A1(\decoded_imm[4] ),
    .A2(_07953_),
    .B1(_07970_),
    .B2(_07971_),
    .X(_01362_));
 sky130_fd_sc_hd__and2_1 _29096_ (.A(\mem_rdata_q[23] ),
    .B(_07850_),
    .X(_07972_));
 sky130_fd_sc_hd__a221o_1 _29097_ (.A1(_07954_),
    .A2(\decoded_imm_uj[3] ),
    .B1(_07929_),
    .B2(\mem_rdata_q[10] ),
    .C1(_07729_),
    .X(_07973_));
 sky130_fd_sc_hd__o22a_1 _29098_ (.A1(\decoded_imm[3] ),
    .A2(_07739_),
    .B1(_07972_),
    .B2(_07973_),
    .X(_01363_));
 sky130_fd_sc_hd__and2_1 _29099_ (.A(\mem_rdata_q[22] ),
    .B(_07850_),
    .X(_07974_));
 sky130_fd_sc_hd__a221o_1 _29100_ (.A1(_06455_),
    .A2(\decoded_imm_uj[2] ),
    .B1(_07929_),
    .B2(\mem_rdata_q[9] ),
    .C1(_07927_),
    .X(_07975_));
 sky130_fd_sc_hd__o22a_1 _29101_ (.A1(\decoded_imm[2] ),
    .A2(_07739_),
    .B1(_07974_),
    .B2(_07975_),
    .X(_01364_));
 sky130_fd_sc_hd__and2_1 _29102_ (.A(\mem_rdata_q[21] ),
    .B(_07850_),
    .X(_07976_));
 sky130_fd_sc_hd__a221o_1 _29103_ (.A1(_06455_),
    .A2(_08546_),
    .B1(_07929_),
    .B2(\mem_rdata_q[8] ),
    .C1(_07927_),
    .X(_07977_));
 sky130_fd_sc_hd__o22a_1 _29104_ (.A1(_08762_),
    .A2(_07739_),
    .B1(_07976_),
    .B2(_07977_),
    .X(_01365_));
 sky130_fd_sc_hd__nor2_1 _29105_ (.A(_08499_),
    .B(_07389_),
    .Y(_01366_));
 sky130_fd_sc_hd__o211ai_2 _29106_ (.A1(_08295_),
    .A2(_08314_),
    .B1(_07679_),
    .C1(_08146_),
    .Y(_07978_));
 sky130_fd_sc_hd__or2_1 _29107_ (.A(_08178_),
    .B(_07978_),
    .X(_07979_));
 sky130_fd_sc_hd__clkbuf_2 _29108_ (.A(_07979_),
    .X(_07980_));
 sky130_fd_sc_hd__and3b_1 _29109_ (.A_N(_07980_),
    .B(_09299_),
    .C(_06578_),
    .X(_07981_));
 sky130_fd_sc_hd__a22o_1 _29110_ (.A1(\latched_rd[3] ),
    .A2(_07980_),
    .B1(_07981_),
    .B2(net444),
    .X(_01367_));
 sky130_fd_sc_hd__a22o_1 _29111_ (.A1(\latched_rd[2] ),
    .A2(_07980_),
    .B1(_07981_),
    .B2(net441),
    .X(_01368_));
 sky130_fd_sc_hd__a22o_1 _29112_ (.A1(\latched_rd[1] ),
    .A2(_07980_),
    .B1(_07981_),
    .B2(net446),
    .X(_01369_));
 sky130_fd_sc_hd__and4bb_1 _29113_ (.A_N(_07323_),
    .B_N(_07978_),
    .C(_06125_),
    .D(_09299_),
    .X(_07982_));
 sky130_fd_sc_hd__a221o_1 _29114_ (.A1(\latched_rd[0] ),
    .A2(_07980_),
    .B1(_07981_),
    .B2(net451),
    .C1(_07982_),
    .X(_01370_));
 sky130_fd_sc_hd__o211a_1 _29115_ (.A1(_06117_),
    .A2(_06405_),
    .B1(_07328_),
    .C1(_08667_),
    .X(_01371_));
 sky130_fd_sc_hd__or2_1 _29116_ (.A(_05268_),
    .B(_05866_),
    .X(_07983_));
 sky130_fd_sc_hd__clkbuf_4 _29117_ (.A(_07983_),
    .X(_07984_));
 sky130_fd_sc_hd__clkbuf_2 _29118_ (.A(_07984_),
    .X(_07985_));
 sky130_fd_sc_hd__mux2_1 _29119_ (.A0(_04988_),
    .A1(\cpuregs[19][0] ),
    .S(_07985_),
    .X(_07986_));
 sky130_fd_sc_hd__clkbuf_1 _29120_ (.A(_07986_),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _29121_ (.A0(_05006_),
    .A1(\cpuregs[19][1] ),
    .S(_07985_),
    .X(_07987_));
 sky130_fd_sc_hd__clkbuf_1 _29122_ (.A(_07987_),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _29123_ (.A0(_05016_),
    .A1(\cpuregs[19][2] ),
    .S(_07985_),
    .X(_07988_));
 sky130_fd_sc_hd__clkbuf_1 _29124_ (.A(_07988_),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _29125_ (.A0(_05023_),
    .A1(\cpuregs[19][3] ),
    .S(_07985_),
    .X(_07989_));
 sky130_fd_sc_hd__clkbuf_1 _29126_ (.A(_07989_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _29127_ (.A0(_05032_),
    .A1(\cpuregs[19][4] ),
    .S(_07985_),
    .X(_07990_));
 sky130_fd_sc_hd__clkbuf_1 _29128_ (.A(_07990_),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _29129_ (.A0(_05041_),
    .A1(\cpuregs[19][5] ),
    .S(_07985_),
    .X(_07991_));
 sky130_fd_sc_hd__clkbuf_1 _29130_ (.A(_07991_),
    .X(_01377_));
 sky130_fd_sc_hd__buf_2 _29131_ (.A(_07984_),
    .X(_07992_));
 sky130_fd_sc_hd__mux2_1 _29132_ (.A0(_05049_),
    .A1(\cpuregs[19][6] ),
    .S(_07992_),
    .X(_07993_));
 sky130_fd_sc_hd__clkbuf_1 _29133_ (.A(_07993_),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _29134_ (.A0(_05060_),
    .A1(\cpuregs[19][7] ),
    .S(_07992_),
    .X(_07994_));
 sky130_fd_sc_hd__clkbuf_1 _29135_ (.A(_07994_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _29136_ (.A0(_05069_),
    .A1(\cpuregs[19][8] ),
    .S(_07992_),
    .X(_07995_));
 sky130_fd_sc_hd__clkbuf_1 _29137_ (.A(_07995_),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_1 _29138_ (.A0(_05076_),
    .A1(\cpuregs[19][9] ),
    .S(_07992_),
    .X(_07996_));
 sky130_fd_sc_hd__clkbuf_1 _29139_ (.A(_07996_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _29140_ (.A0(_05085_),
    .A1(\cpuregs[19][10] ),
    .S(_07992_),
    .X(_07997_));
 sky130_fd_sc_hd__clkbuf_1 _29141_ (.A(_07997_),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _29142_ (.A0(_05095_),
    .A1(\cpuregs[19][11] ),
    .S(_07992_),
    .X(_07998_));
 sky130_fd_sc_hd__clkbuf_1 _29143_ (.A(_07998_),
    .X(_01383_));
 sky130_fd_sc_hd__clkbuf_2 _29144_ (.A(_07984_),
    .X(_07999_));
 sky130_fd_sc_hd__mux2_1 _29145_ (.A0(_05102_),
    .A1(\cpuregs[19][12] ),
    .S(_07999_),
    .X(_08000_));
 sky130_fd_sc_hd__clkbuf_1 _29146_ (.A(_08000_),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_1 _29147_ (.A0(_05113_),
    .A1(\cpuregs[19][13] ),
    .S(_07999_),
    .X(_08001_));
 sky130_fd_sc_hd__clkbuf_1 _29148_ (.A(_08001_),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _29149_ (.A0(_05121_),
    .A1(\cpuregs[19][14] ),
    .S(_07999_),
    .X(_08002_));
 sky130_fd_sc_hd__clkbuf_1 _29150_ (.A(_08002_),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _29151_ (.A0(_05129_),
    .A1(\cpuregs[19][15] ),
    .S(_07999_),
    .X(_08003_));
 sky130_fd_sc_hd__clkbuf_1 _29152_ (.A(_08003_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _29153_ (.A0(_05138_),
    .A1(\cpuregs[19][16] ),
    .S(_07999_),
    .X(_08004_));
 sky130_fd_sc_hd__clkbuf_1 _29154_ (.A(_08004_),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _29155_ (.A0(_05146_),
    .A1(\cpuregs[19][17] ),
    .S(_07999_),
    .X(_08005_));
 sky130_fd_sc_hd__clkbuf_1 _29156_ (.A(_08005_),
    .X(_01389_));
 sky130_fd_sc_hd__clkbuf_2 _29157_ (.A(_07984_),
    .X(_08006_));
 sky130_fd_sc_hd__mux2_1 _29158_ (.A0(_05154_),
    .A1(\cpuregs[19][18] ),
    .S(_08006_),
    .X(_08007_));
 sky130_fd_sc_hd__clkbuf_1 _29159_ (.A(_08007_),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_1 _29160_ (.A0(_05165_),
    .A1(\cpuregs[19][19] ),
    .S(_08006_),
    .X(_08008_));
 sky130_fd_sc_hd__clkbuf_1 _29161_ (.A(_08008_),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _29162_ (.A0(_05173_),
    .A1(\cpuregs[19][20] ),
    .S(_08006_),
    .X(_08009_));
 sky130_fd_sc_hd__clkbuf_1 _29163_ (.A(_08009_),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _29164_ (.A0(_05182_),
    .A1(\cpuregs[19][21] ),
    .S(_08006_),
    .X(_08010_));
 sky130_fd_sc_hd__clkbuf_1 _29165_ (.A(_08010_),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _29166_ (.A0(_05191_),
    .A1(\cpuregs[19][22] ),
    .S(_08006_),
    .X(_08011_));
 sky130_fd_sc_hd__clkbuf_1 _29167_ (.A(_08011_),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _29168_ (.A0(_05199_),
    .A1(\cpuregs[19][23] ),
    .S(_08006_),
    .X(_08012_));
 sky130_fd_sc_hd__clkbuf_1 _29169_ (.A(_08012_),
    .X(_01395_));
 sky130_fd_sc_hd__buf_2 _29170_ (.A(_07983_),
    .X(_08013_));
 sky130_fd_sc_hd__mux2_1 _29171_ (.A0(_05206_),
    .A1(\cpuregs[19][24] ),
    .S(_08013_),
    .X(_08014_));
 sky130_fd_sc_hd__clkbuf_1 _29172_ (.A(_08014_),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _29173_ (.A0(_05217_),
    .A1(\cpuregs[19][25] ),
    .S(_08013_),
    .X(_08015_));
 sky130_fd_sc_hd__clkbuf_1 _29174_ (.A(_08015_),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _29175_ (.A0(_05225_),
    .A1(\cpuregs[19][26] ),
    .S(_08013_),
    .X(_08016_));
 sky130_fd_sc_hd__clkbuf_1 _29176_ (.A(_08016_),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _29177_ (.A0(_05232_),
    .A1(\cpuregs[19][27] ),
    .S(_08013_),
    .X(_08017_));
 sky130_fd_sc_hd__clkbuf_1 _29178_ (.A(_08017_),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _29179_ (.A0(_05240_),
    .A1(\cpuregs[19][28] ),
    .S(_08013_),
    .X(_08018_));
 sky130_fd_sc_hd__clkbuf_1 _29180_ (.A(_08018_),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _29181_ (.A0(_05248_),
    .A1(\cpuregs[19][29] ),
    .S(_08013_),
    .X(_08019_));
 sky130_fd_sc_hd__clkbuf_1 _29182_ (.A(_08019_),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _29183_ (.A0(_05256_),
    .A1(\cpuregs[19][30] ),
    .S(_07984_),
    .X(_08020_));
 sky130_fd_sc_hd__clkbuf_1 _29184_ (.A(_08020_),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _29185_ (.A0(_05263_),
    .A1(\cpuregs[19][31] ),
    .S(_07984_),
    .X(_08021_));
 sky130_fd_sc_hd__clkbuf_1 _29186_ (.A(_08021_),
    .X(_01403_));
 sky130_fd_sc_hd__o21a_1 _29187_ (.A1(\decoded_rd[4] ),
    .A2(_06620_),
    .B1(_09299_),
    .X(_08022_));
 sky130_fd_sc_hd__o21ba_1 _29188_ (.A1(_06125_),
    .A2(instr_setq),
    .B1_N(_07978_),
    .X(_08023_));
 sky130_fd_sc_hd__o22a_1 _29189_ (.A1(_07980_),
    .A2(_08022_),
    .B1(_08023_),
    .B2(\latched_rd[4] ),
    .X(_01404_));
 sky130_fd_sc_hd__o2bb2a_1 _29190_ (.A1_N(_05548_),
    .A2_N(_07832_),
    .B1(\decoded_rs1[4] ),
    .B2(_05538_),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _29191_ (.A0(net119),
    .A1(net150),
    .S(_05748_),
    .X(_08024_));
 sky130_fd_sc_hd__clkbuf_1 _29192_ (.A(_08024_),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _29193_ (.A0(net122),
    .A1(net153),
    .S(_05748_),
    .X(_08025_));
 sky130_fd_sc_hd__clkbuf_1 _29194_ (.A(_08025_),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _29195_ (.A0(net123),
    .A1(net154),
    .S(_05748_),
    .X(_08026_));
 sky130_fd_sc_hd__clkbuf_1 _29196_ (.A(_08026_),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _29197_ (.A0(net124),
    .A1(net155),
    .S(_05748_),
    .X(_08027_));
 sky130_fd_sc_hd__clkbuf_1 _29198_ (.A(_08027_),
    .X(_01409_));
 sky130_fd_sc_hd__clkbuf_2 _29199_ (.A(_05747_),
    .X(_08028_));
 sky130_fd_sc_hd__mux2_1 _29200_ (.A0(net125),
    .A1(net156),
    .S(_08028_),
    .X(_08029_));
 sky130_fd_sc_hd__clkbuf_1 _29201_ (.A(_08029_),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _29202_ (.A0(net126),
    .A1(net157),
    .S(_08028_),
    .X(_08030_));
 sky130_fd_sc_hd__clkbuf_1 _29203_ (.A(_08030_),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _29204_ (.A0(net127),
    .A1(net158),
    .S(_08028_),
    .X(_08031_));
 sky130_fd_sc_hd__clkbuf_1 _29205_ (.A(_08031_),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _29206_ (.A0(net128),
    .A1(net159),
    .S(_08028_),
    .X(_08032_));
 sky130_fd_sc_hd__clkbuf_1 _29207_ (.A(_08032_),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_1 _29208_ (.A0(net99),
    .A1(net130),
    .S(_08028_),
    .X(_08033_));
 sky130_fd_sc_hd__clkbuf_1 _29209_ (.A(_08033_),
    .X(_01414_));
 sky130_fd_sc_hd__mux2_1 _29210_ (.A0(net100),
    .A1(net131),
    .S(_08028_),
    .X(_08034_));
 sky130_fd_sc_hd__clkbuf_1 _29211_ (.A(_08034_),
    .X(_01415_));
 sky130_fd_sc_hd__clkbuf_2 _29212_ (.A(_05747_),
    .X(_08035_));
 sky130_fd_sc_hd__mux2_1 _29213_ (.A0(net101),
    .A1(net132),
    .S(_08035_),
    .X(_08036_));
 sky130_fd_sc_hd__clkbuf_1 _29214_ (.A(_08036_),
    .X(_01416_));
 sky130_fd_sc_hd__mux2_1 _29215_ (.A0(net102),
    .A1(net133),
    .S(_08035_),
    .X(_08037_));
 sky130_fd_sc_hd__clkbuf_1 _29216_ (.A(_08037_),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _29217_ (.A0(net103),
    .A1(net134),
    .S(_08035_),
    .X(_08038_));
 sky130_fd_sc_hd__clkbuf_1 _29218_ (.A(_08038_),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _29219_ (.A0(net104),
    .A1(net135),
    .S(_08035_),
    .X(_08039_));
 sky130_fd_sc_hd__clkbuf_1 _29220_ (.A(_08039_),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _29221_ (.A0(net105),
    .A1(net136),
    .S(_08035_),
    .X(_08040_));
 sky130_fd_sc_hd__clkbuf_1 _29222_ (.A(_08040_),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _29223_ (.A0(net106),
    .A1(net137),
    .S(_08035_),
    .X(_08041_));
 sky130_fd_sc_hd__clkbuf_1 _29224_ (.A(_08041_),
    .X(_01421_));
 sky130_fd_sc_hd__buf_2 _29225_ (.A(_05747_),
    .X(_08042_));
 sky130_fd_sc_hd__mux2_1 _29226_ (.A0(net107),
    .A1(net138),
    .S(_08042_),
    .X(_08043_));
 sky130_fd_sc_hd__clkbuf_1 _29227_ (.A(_08043_),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _29228_ (.A0(net108),
    .A1(net139),
    .S(_08042_),
    .X(_08044_));
 sky130_fd_sc_hd__clkbuf_1 _29229_ (.A(_08044_),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_1 _29230_ (.A0(net109),
    .A1(net140),
    .S(_08042_),
    .X(_08045_));
 sky130_fd_sc_hd__clkbuf_1 _29231_ (.A(_08045_),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _29232_ (.A0(net110),
    .A1(net141),
    .S(_08042_),
    .X(_08046_));
 sky130_fd_sc_hd__clkbuf_1 _29233_ (.A(_08046_),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _29234_ (.A0(net111),
    .A1(net142),
    .S(_08042_),
    .X(_08047_));
 sky130_fd_sc_hd__clkbuf_1 _29235_ (.A(_08047_),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_1 _29236_ (.A0(net112),
    .A1(net143),
    .S(_08042_),
    .X(_08048_));
 sky130_fd_sc_hd__clkbuf_1 _29237_ (.A(_08048_),
    .X(_01427_));
 sky130_fd_sc_hd__buf_2 _29238_ (.A(_05746_),
    .X(_08049_));
 sky130_fd_sc_hd__mux2_1 _29239_ (.A0(net113),
    .A1(net144),
    .S(_08049_),
    .X(_08050_));
 sky130_fd_sc_hd__clkbuf_1 _29240_ (.A(_08050_),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_1 _29241_ (.A0(net114),
    .A1(net145),
    .S(_08049_),
    .X(_08051_));
 sky130_fd_sc_hd__clkbuf_1 _29242_ (.A(_08051_),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _29243_ (.A0(net115),
    .A1(net146),
    .S(_08049_),
    .X(_08052_));
 sky130_fd_sc_hd__clkbuf_1 _29244_ (.A(_08052_),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _29245_ (.A0(net116),
    .A1(net147),
    .S(_08049_),
    .X(_08053_));
 sky130_fd_sc_hd__clkbuf_1 _29246_ (.A(_08053_),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_1 _29247_ (.A0(net117),
    .A1(net148),
    .S(_08049_),
    .X(_08054_));
 sky130_fd_sc_hd__clkbuf_1 _29248_ (.A(_08054_),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _29249_ (.A0(net118),
    .A1(net149),
    .S(_08049_),
    .X(_08055_));
 sky130_fd_sc_hd__clkbuf_1 _29250_ (.A(_08055_),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _29251_ (.A0(net120),
    .A1(net151),
    .S(_05747_),
    .X(_08056_));
 sky130_fd_sc_hd__clkbuf_1 _29252_ (.A(_08056_),
    .X(_01434_));
 sky130_fd_sc_hd__mux2_1 _29253_ (.A0(net121),
    .A1(net152),
    .S(_05747_),
    .X(_08057_));
 sky130_fd_sc_hd__clkbuf_1 _29254_ (.A(_08057_),
    .X(_01435_));
 sky130_fd_sc_hd__nor2_1 _29255_ (.A(_05340_),
    .B(_05468_),
    .Y(_08058_));
 sky130_fd_sc_hd__clkbuf_4 _29256_ (.A(_08058_),
    .X(_08059_));
 sky130_fd_sc_hd__buf_2 _29257_ (.A(_08059_),
    .X(_08060_));
 sky130_fd_sc_hd__mux2_1 _29258_ (.A0(\cpuregs[9][0] ),
    .A1(_05665_),
    .S(_08060_),
    .X(_08061_));
 sky130_fd_sc_hd__clkbuf_1 _29259_ (.A(_08061_),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _29260_ (.A0(\cpuregs[9][1] ),
    .A1(_05671_),
    .S(_08060_),
    .X(_08062_));
 sky130_fd_sc_hd__clkbuf_1 _29261_ (.A(_08062_),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _29262_ (.A0(\cpuregs[9][2] ),
    .A1(_05673_),
    .S(_08060_),
    .X(_08063_));
 sky130_fd_sc_hd__clkbuf_1 _29263_ (.A(_08063_),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _29264_ (.A0(\cpuregs[9][3] ),
    .A1(_05675_),
    .S(_08060_),
    .X(_08064_));
 sky130_fd_sc_hd__clkbuf_1 _29265_ (.A(_08064_),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _29266_ (.A0(\cpuregs[9][4] ),
    .A1(_05677_),
    .S(_08060_),
    .X(_08065_));
 sky130_fd_sc_hd__clkbuf_1 _29267_ (.A(_08065_),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_1 _29268_ (.A0(\cpuregs[9][5] ),
    .A1(_05679_),
    .S(_08060_),
    .X(_08066_));
 sky130_fd_sc_hd__clkbuf_1 _29269_ (.A(_08066_),
    .X(_01441_));
 sky130_fd_sc_hd__buf_2 _29270_ (.A(_08059_),
    .X(_08067_));
 sky130_fd_sc_hd__mux2_1 _29271_ (.A0(\cpuregs[9][6] ),
    .A1(_05681_),
    .S(_08067_),
    .X(_08068_));
 sky130_fd_sc_hd__clkbuf_1 _29272_ (.A(_08068_),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _29273_ (.A0(\cpuregs[9][7] ),
    .A1(_05684_),
    .S(_08067_),
    .X(_08069_));
 sky130_fd_sc_hd__clkbuf_1 _29274_ (.A(_08069_),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_1 _29275_ (.A0(\cpuregs[9][8] ),
    .A1(_05686_),
    .S(_08067_),
    .X(_08070_));
 sky130_fd_sc_hd__clkbuf_1 _29276_ (.A(_08070_),
    .X(_01444_));
 sky130_fd_sc_hd__mux2_1 _29277_ (.A0(\cpuregs[9][9] ),
    .A1(_05688_),
    .S(_08067_),
    .X(_08071_));
 sky130_fd_sc_hd__clkbuf_1 _29278_ (.A(_08071_),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _29279_ (.A0(\cpuregs[9][10] ),
    .A1(_05690_),
    .S(_08067_),
    .X(_08072_));
 sky130_fd_sc_hd__clkbuf_1 _29280_ (.A(_08072_),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_1 _29281_ (.A0(\cpuregs[9][11] ),
    .A1(_05692_),
    .S(_08067_),
    .X(_08073_));
 sky130_fd_sc_hd__clkbuf_1 _29282_ (.A(_08073_),
    .X(_01447_));
 sky130_fd_sc_hd__clkbuf_4 _29283_ (.A(_08059_),
    .X(_08074_));
 sky130_fd_sc_hd__mux2_1 _29284_ (.A0(\cpuregs[9][12] ),
    .A1(_05694_),
    .S(_08074_),
    .X(_08075_));
 sky130_fd_sc_hd__clkbuf_1 _29285_ (.A(_08075_),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _29286_ (.A0(\cpuregs[9][13] ),
    .A1(_05697_),
    .S(_08074_),
    .X(_08076_));
 sky130_fd_sc_hd__clkbuf_1 _29287_ (.A(_08076_),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _29288_ (.A0(\cpuregs[9][14] ),
    .A1(_05699_),
    .S(_08074_),
    .X(_08077_));
 sky130_fd_sc_hd__clkbuf_1 _29289_ (.A(_08077_),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _29290_ (.A0(\cpuregs[9][15] ),
    .A1(_05701_),
    .S(_08074_),
    .X(_08078_));
 sky130_fd_sc_hd__clkbuf_1 _29291_ (.A(_08078_),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _29292_ (.A0(\cpuregs[9][16] ),
    .A1(_05703_),
    .S(_08074_),
    .X(_08079_));
 sky130_fd_sc_hd__clkbuf_1 _29293_ (.A(_08079_),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_1 _29294_ (.A0(\cpuregs[9][17] ),
    .A1(_05705_),
    .S(_08074_),
    .X(_08080_));
 sky130_fd_sc_hd__clkbuf_1 _29295_ (.A(_08080_),
    .X(_01453_));
 sky130_fd_sc_hd__buf_2 _29296_ (.A(_08059_),
    .X(_08081_));
 sky130_fd_sc_hd__mux2_1 _29297_ (.A0(\cpuregs[9][18] ),
    .A1(_05707_),
    .S(_08081_),
    .X(_08082_));
 sky130_fd_sc_hd__clkbuf_1 _29298_ (.A(_08082_),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _29299_ (.A0(\cpuregs[9][19] ),
    .A1(_05710_),
    .S(_08081_),
    .X(_08083_));
 sky130_fd_sc_hd__clkbuf_1 _29300_ (.A(_08083_),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _29301_ (.A0(\cpuregs[9][20] ),
    .A1(_05712_),
    .S(_08081_),
    .X(_08084_));
 sky130_fd_sc_hd__clkbuf_1 _29302_ (.A(_08084_),
    .X(_01456_));
 sky130_fd_sc_hd__mux2_1 _29303_ (.A0(\cpuregs[9][21] ),
    .A1(_05714_),
    .S(_08081_),
    .X(_08085_));
 sky130_fd_sc_hd__clkbuf_1 _29304_ (.A(_08085_),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _29305_ (.A0(\cpuregs[9][22] ),
    .A1(_05716_),
    .S(_08081_),
    .X(_08086_));
 sky130_fd_sc_hd__clkbuf_1 _29306_ (.A(_08086_),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _29307_ (.A0(\cpuregs[9][23] ),
    .A1(_05718_),
    .S(_08081_),
    .X(_08087_));
 sky130_fd_sc_hd__clkbuf_1 _29308_ (.A(_08087_),
    .X(_01459_));
 sky130_fd_sc_hd__clkbuf_4 _29309_ (.A(_08058_),
    .X(_08088_));
 sky130_fd_sc_hd__mux2_1 _29310_ (.A0(\cpuregs[9][24] ),
    .A1(_05720_),
    .S(_08088_),
    .X(_08089_));
 sky130_fd_sc_hd__clkbuf_1 _29311_ (.A(_08089_),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _29312_ (.A0(\cpuregs[9][25] ),
    .A1(_05723_),
    .S(_08088_),
    .X(_08090_));
 sky130_fd_sc_hd__clkbuf_1 _29313_ (.A(_08090_),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _29314_ (.A0(\cpuregs[9][26] ),
    .A1(_05725_),
    .S(_08088_),
    .X(_08091_));
 sky130_fd_sc_hd__clkbuf_1 _29315_ (.A(_08091_),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_1 _29316_ (.A0(\cpuregs[9][27] ),
    .A1(_05727_),
    .S(_08088_),
    .X(_08092_));
 sky130_fd_sc_hd__clkbuf_1 _29317_ (.A(_08092_),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _29318_ (.A0(\cpuregs[9][28] ),
    .A1(_05729_),
    .S(_08088_),
    .X(_08093_));
 sky130_fd_sc_hd__clkbuf_1 _29319_ (.A(_08093_),
    .X(_01464_));
 sky130_fd_sc_hd__mux2_1 _29320_ (.A0(\cpuregs[9][29] ),
    .A1(_05731_),
    .S(_08088_),
    .X(_08094_));
 sky130_fd_sc_hd__clkbuf_1 _29321_ (.A(_08094_),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _29322_ (.A0(\cpuregs[9][30] ),
    .A1(_05733_),
    .S(_08059_),
    .X(_08095_));
 sky130_fd_sc_hd__clkbuf_1 _29323_ (.A(_08095_),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _29324_ (.A0(\cpuregs[9][31] ),
    .A1(_05735_),
    .S(_08059_),
    .X(_08096_));
 sky130_fd_sc_hd__clkbuf_1 _29325_ (.A(_08096_),
    .X(_01467_));
 sky130_fd_sc_hd__nor2_1 _29326_ (.A(_05269_),
    .B(_05340_),
    .Y(_08097_));
 sky130_fd_sc_hd__buf_4 _29327_ (.A(_08097_),
    .X(_08098_));
 sky130_fd_sc_hd__buf_2 _29328_ (.A(_08098_),
    .X(_08099_));
 sky130_fd_sc_hd__mux2_1 _29329_ (.A0(\cpuregs[1][0] ),
    .A1(_04987_),
    .S(_08099_),
    .X(_08100_));
 sky130_fd_sc_hd__clkbuf_1 _29330_ (.A(_08100_),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _29331_ (.A0(\cpuregs[1][1] ),
    .A1(_05005_),
    .S(_08099_),
    .X(_08101_));
 sky130_fd_sc_hd__clkbuf_1 _29332_ (.A(_08101_),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _29333_ (.A0(\cpuregs[1][2] ),
    .A1(_05015_),
    .S(_08099_),
    .X(_08102_));
 sky130_fd_sc_hd__clkbuf_1 _29334_ (.A(_08102_),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _29335_ (.A0(\cpuregs[1][3] ),
    .A1(_05022_),
    .S(_08099_),
    .X(_08103_));
 sky130_fd_sc_hd__clkbuf_1 _29336_ (.A(_08103_),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _29337_ (.A0(\cpuregs[1][4] ),
    .A1(_05031_),
    .S(_08099_),
    .X(_08104_));
 sky130_fd_sc_hd__clkbuf_1 _29338_ (.A(_08104_),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _29339_ (.A0(\cpuregs[1][5] ),
    .A1(_05040_),
    .S(_08099_),
    .X(_08105_));
 sky130_fd_sc_hd__clkbuf_1 _29340_ (.A(_08105_),
    .X(_01473_));
 sky130_fd_sc_hd__clkbuf_4 _29341_ (.A(_08098_),
    .X(_08106_));
 sky130_fd_sc_hd__mux2_1 _29342_ (.A0(\cpuregs[1][6] ),
    .A1(_05048_),
    .S(_08106_),
    .X(_08107_));
 sky130_fd_sc_hd__clkbuf_1 _29343_ (.A(_08107_),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_1 _29344_ (.A0(\cpuregs[1][7] ),
    .A1(_05059_),
    .S(_08106_),
    .X(_08108_));
 sky130_fd_sc_hd__clkbuf_1 _29345_ (.A(_08108_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _29346_ (.A0(\cpuregs[1][8] ),
    .A1(_05068_),
    .S(_08106_),
    .X(_08109_));
 sky130_fd_sc_hd__clkbuf_1 _29347_ (.A(_08109_),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _29348_ (.A0(\cpuregs[1][9] ),
    .A1(_05075_),
    .S(_08106_),
    .X(_08110_));
 sky130_fd_sc_hd__clkbuf_1 _29349_ (.A(_08110_),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _29350_ (.A0(\cpuregs[1][10] ),
    .A1(_05084_),
    .S(_08106_),
    .X(_08111_));
 sky130_fd_sc_hd__clkbuf_1 _29351_ (.A(_08111_),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _29352_ (.A0(\cpuregs[1][11] ),
    .A1(_05094_),
    .S(_08106_),
    .X(_08112_));
 sky130_fd_sc_hd__clkbuf_1 _29353_ (.A(_08112_),
    .X(_01479_));
 sky130_fd_sc_hd__clkbuf_4 _29354_ (.A(_08098_),
    .X(_08113_));
 sky130_fd_sc_hd__mux2_1 _29355_ (.A0(\cpuregs[1][12] ),
    .A1(_05101_),
    .S(_08113_),
    .X(_08114_));
 sky130_fd_sc_hd__clkbuf_1 _29356_ (.A(_08114_),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _29357_ (.A0(\cpuregs[1][13] ),
    .A1(_05112_),
    .S(_08113_),
    .X(_08115_));
 sky130_fd_sc_hd__clkbuf_1 _29358_ (.A(_08115_),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _29359_ (.A0(\cpuregs[1][14] ),
    .A1(_05120_),
    .S(_08113_),
    .X(_08116_));
 sky130_fd_sc_hd__clkbuf_1 _29360_ (.A(_08116_),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _29361_ (.A0(\cpuregs[1][15] ),
    .A1(_05128_),
    .S(_08113_),
    .X(_08117_));
 sky130_fd_sc_hd__clkbuf_1 _29362_ (.A(_08117_),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _29363_ (.A0(\cpuregs[1][16] ),
    .A1(_05137_),
    .S(_08113_),
    .X(_08118_));
 sky130_fd_sc_hd__clkbuf_1 _29364_ (.A(_08118_),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_1 _29365_ (.A0(\cpuregs[1][17] ),
    .A1(_05145_),
    .S(_08113_),
    .X(_08119_));
 sky130_fd_sc_hd__clkbuf_1 _29366_ (.A(_08119_),
    .X(_01485_));
 sky130_fd_sc_hd__buf_2 _29367_ (.A(_08098_),
    .X(_08120_));
 sky130_fd_sc_hd__mux2_1 _29368_ (.A0(\cpuregs[1][18] ),
    .A1(_05153_),
    .S(_08120_),
    .X(_08121_));
 sky130_fd_sc_hd__clkbuf_1 _29369_ (.A(_08121_),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _29370_ (.A0(\cpuregs[1][19] ),
    .A1(_05164_),
    .S(_08120_),
    .X(_08122_));
 sky130_fd_sc_hd__clkbuf_1 _29371_ (.A(_08122_),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _29372_ (.A0(\cpuregs[1][20] ),
    .A1(_05172_),
    .S(_08120_),
    .X(_08123_));
 sky130_fd_sc_hd__clkbuf_1 _29373_ (.A(_08123_),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _29374_ (.A0(\cpuregs[1][21] ),
    .A1(_05181_),
    .S(_08120_),
    .X(_08124_));
 sky130_fd_sc_hd__clkbuf_1 _29375_ (.A(_08124_),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _29376_ (.A0(\cpuregs[1][22] ),
    .A1(_05190_),
    .S(_08120_),
    .X(_08125_));
 sky130_fd_sc_hd__clkbuf_1 _29377_ (.A(_08125_),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _29378_ (.A0(\cpuregs[1][23] ),
    .A1(_05198_),
    .S(_08120_),
    .X(_08126_));
 sky130_fd_sc_hd__clkbuf_1 _29379_ (.A(_08126_),
    .X(_01491_));
 sky130_fd_sc_hd__clkbuf_4 _29380_ (.A(_08097_),
    .X(_08127_));
 sky130_fd_sc_hd__mux2_1 _29381_ (.A0(\cpuregs[1][24] ),
    .A1(_05205_),
    .S(_08127_),
    .X(_08128_));
 sky130_fd_sc_hd__clkbuf_1 _29382_ (.A(_08128_),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _29383_ (.A0(\cpuregs[1][25] ),
    .A1(_05216_),
    .S(_08127_),
    .X(_08129_));
 sky130_fd_sc_hd__clkbuf_1 _29384_ (.A(_08129_),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _29385_ (.A0(\cpuregs[1][26] ),
    .A1(_05224_),
    .S(_08127_),
    .X(_08130_));
 sky130_fd_sc_hd__clkbuf_1 _29386_ (.A(_08130_),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _29387_ (.A0(\cpuregs[1][27] ),
    .A1(_05231_),
    .S(_08127_),
    .X(_08131_));
 sky130_fd_sc_hd__clkbuf_1 _29388_ (.A(_08131_),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _29389_ (.A0(\cpuregs[1][28] ),
    .A1(_05239_),
    .S(_08127_),
    .X(_08132_));
 sky130_fd_sc_hd__clkbuf_1 _29390_ (.A(_08132_),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _29391_ (.A0(\cpuregs[1][29] ),
    .A1(_05247_),
    .S(_08127_),
    .X(_08133_));
 sky130_fd_sc_hd__clkbuf_1 _29392_ (.A(_08133_),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _29393_ (.A0(\cpuregs[1][30] ),
    .A1(_05255_),
    .S(_08098_),
    .X(_08134_));
 sky130_fd_sc_hd__clkbuf_1 _29394_ (.A(_08134_),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _29395_ (.A0(\cpuregs[1][31] ),
    .A1(_05262_),
    .S(_08098_),
    .X(_08135_));
 sky130_fd_sc_hd__clkbuf_1 _29396_ (.A(_08135_),
    .X(_01499_));
 sky130_fd_sc_hd__dfxtp_1 _29397_ (.CLK(clknet_leaf_186_clk),
    .D(_00114_),
    .Q(\cpuregs[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29398_ (.CLK(clknet_leaf_181_clk),
    .D(_00115_),
    .Q(\cpuregs[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29399_ (.CLK(clknet_leaf_180_clk),
    .D(_00116_),
    .Q(\cpuregs[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29400_ (.CLK(clknet_leaf_180_clk),
    .D(_00117_),
    .Q(\cpuregs[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29401_ (.CLK(clknet_leaf_179_clk),
    .D(_00118_),
    .Q(\cpuregs[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29402_ (.CLK(clknet_leaf_184_clk),
    .D(_00119_),
    .Q(\cpuregs[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29403_ (.CLK(clknet_leaf_184_clk),
    .D(_00120_),
    .Q(\cpuregs[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29404_ (.CLK(clknet_leaf_191_clk),
    .D(_00121_),
    .Q(\cpuregs[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29405_ (.CLK(clknet_leaf_154_clk),
    .D(_00122_),
    .Q(\cpuregs[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29406_ (.CLK(clknet_leaf_156_clk),
    .D(_00123_),
    .Q(\cpuregs[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29407_ (.CLK(clknet_leaf_189_clk),
    .D(_00124_),
    .Q(\cpuregs[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29408_ (.CLK(clknet_leaf_183_clk),
    .D(_00125_),
    .Q(\cpuregs[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29409_ (.CLK(clknet_leaf_123_clk),
    .D(_00126_),
    .Q(\cpuregs[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29410_ (.CLK(clknet_leaf_101_clk),
    .D(_00127_),
    .Q(\cpuregs[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29411_ (.CLK(clknet_leaf_100_clk),
    .D(_00128_),
    .Q(\cpuregs[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29412_ (.CLK(clknet_leaf_140_clk),
    .D(_00129_),
    .Q(\cpuregs[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29413_ (.CLK(clknet_leaf_124_clk),
    .D(_00130_),
    .Q(\cpuregs[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29414_ (.CLK(clknet_leaf_121_clk),
    .D(_00131_),
    .Q(\cpuregs[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29415_ (.CLK(clknet_leaf_155_clk),
    .D(_00132_),
    .Q(\cpuregs[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29416_ (.CLK(clknet_leaf_159_clk),
    .D(_00133_),
    .Q(\cpuregs[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29417_ (.CLK(clknet_leaf_155_clk),
    .D(_00134_),
    .Q(\cpuregs[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29418_ (.CLK(clknet_leaf_159_clk),
    .D(_00135_),
    .Q(\cpuregs[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29419_ (.CLK(clknet_leaf_155_clk),
    .D(_00136_),
    .Q(\cpuregs[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29420_ (.CLK(clknet_leaf_155_clk),
    .D(_00137_),
    .Q(\cpuregs[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29421_ (.CLK(clknet_leaf_129_clk),
    .D(_00138_),
    .Q(\cpuregs[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29422_ (.CLK(clknet_leaf_130_clk),
    .D(_00139_),
    .Q(\cpuregs[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29423_ (.CLK(clknet_leaf_119_clk),
    .D(_00140_),
    .Q(\cpuregs[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29424_ (.CLK(clknet_leaf_118_clk),
    .D(_00141_),
    .Q(\cpuregs[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29425_ (.CLK(clknet_leaf_126_clk),
    .D(_00142_),
    .Q(\cpuregs[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29426_ (.CLK(clknet_leaf_127_clk),
    .D(_00143_),
    .Q(\cpuregs[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29427_ (.CLK(clknet_leaf_138_clk),
    .D(_00144_),
    .Q(\cpuregs[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29428_ (.CLK(clknet_leaf_145_clk),
    .D(_00145_),
    .Q(\cpuregs[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29429_ (.CLK(clknet_leaf_159_clk),
    .D(_00146_),
    .Q(\cpuregs[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29430_ (.CLK(clknet_leaf_171_clk),
    .D(_00147_),
    .Q(\cpuregs[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29431_ (.CLK(clknet_leaf_171_clk),
    .D(_00148_),
    .Q(\cpuregs[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29432_ (.CLK(clknet_leaf_169_clk),
    .D(_00149_),
    .Q(\cpuregs[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29433_ (.CLK(clknet_leaf_170_clk),
    .D(_00150_),
    .Q(\cpuregs[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29434_ (.CLK(clknet_leaf_169_clk),
    .D(_00151_),
    .Q(\cpuregs[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29435_ (.CLK(clknet_leaf_184_clk),
    .D(_00152_),
    .Q(\cpuregs[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29436_ (.CLK(clknet_leaf_193_clk),
    .D(_00153_),
    .Q(\cpuregs[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29437_ (.CLK(clknet_leaf_192_clk),
    .D(_00154_),
    .Q(\cpuregs[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29438_ (.CLK(clknet_leaf_192_clk),
    .D(_00155_),
    .Q(\cpuregs[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29439_ (.CLK(clknet_leaf_189_clk),
    .D(_00156_),
    .Q(\cpuregs[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29440_ (.CLK(clknet_leaf_188_clk),
    .D(_00157_),
    .Q(\cpuregs[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29441_ (.CLK(clknet_leaf_135_clk),
    .D(_00158_),
    .Q(\cpuregs[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29442_ (.CLK(clknet_leaf_123_clk),
    .D(_00159_),
    .Q(\cpuregs[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29443_ (.CLK(clknet_leaf_164_clk),
    .D(_00160_),
    .Q(\cpuregs[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29444_ (.CLK(clknet_leaf_141_clk),
    .D(_00161_),
    .Q(\cpuregs[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29445_ (.CLK(clknet_leaf_134_clk),
    .D(_00162_),
    .Q(\cpuregs[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29446_ (.CLK(clknet_leaf_124_clk),
    .D(_00163_),
    .Q(\cpuregs[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29447_ (.CLK(clknet_leaf_144_clk),
    .D(_00164_),
    .Q(\cpuregs[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29448_ (.CLK(clknet_leaf_148_clk),
    .D(_00165_),
    .Q(\cpuregs[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29449_ (.CLK(clknet_leaf_149_clk),
    .D(_00166_),
    .Q(\cpuregs[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29450_ (.CLK(clknet_leaf_147_clk),
    .D(_00167_),
    .Q(\cpuregs[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29451_ (.CLK(clknet_leaf_147_clk),
    .D(_00168_),
    .Q(\cpuregs[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29452_ (.CLK(clknet_leaf_148_clk),
    .D(_00169_),
    .Q(\cpuregs[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29453_ (.CLK(clknet_leaf_129_clk),
    .D(_00170_),
    .Q(\cpuregs[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29454_ (.CLK(clknet_leaf_130_clk),
    .D(_00171_),
    .Q(\cpuregs[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29455_ (.CLK(clknet_leaf_117_clk),
    .D(_00172_),
    .Q(\cpuregs[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29456_ (.CLK(clknet_leaf_118_clk),
    .D(_00173_),
    .Q(\cpuregs[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29457_ (.CLK(clknet_leaf_125_clk),
    .D(_00174_),
    .Q(\cpuregs[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29458_ (.CLK(clknet_leaf_117_clk),
    .D(_00175_),
    .Q(\cpuregs[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29459_ (.CLK(clknet_leaf_134_clk),
    .D(_00176_),
    .Q(\cpuregs[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29460_ (.CLK(clknet_leaf_146_clk),
    .D(_00177_),
    .Q(\cpuregs[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29461_ (.CLK(clknet_leaf_204_clk),
    .D(_00050_),
    .Q(\genblk1.pcpi_mul.rd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _29462_ (.CLK(clknet_leaf_204_clk),
    .D(_00051_),
    .Q(\genblk1.pcpi_mul.rd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _29463_ (.CLK(clknet_leaf_204_clk),
    .D(_00052_),
    .Q(\genblk1.pcpi_mul.rd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _29464_ (.CLK(clknet_leaf_205_clk),
    .D(_00053_),
    .Q(\genblk1.pcpi_mul.rd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _29465_ (.CLK(clknet_leaf_201_clk),
    .D(_00054_),
    .Q(\genblk1.pcpi_mul.rd[4] ));
 sky130_fd_sc_hd__dfxtp_1 _29466_ (.CLK(clknet_leaf_205_clk),
    .D(_00055_),
    .Q(\genblk1.pcpi_mul.rd[5] ));
 sky130_fd_sc_hd__dfxtp_1 _29467_ (.CLK(clknet_leaf_205_clk),
    .D(_00110_),
    .Q(\genblk1.pcpi_mul.rd[6] ));
 sky130_fd_sc_hd__dfxtp_1 _29468_ (.CLK(clknet_leaf_203_clk),
    .D(_00111_),
    .Q(\genblk1.pcpi_mul.rd[7] ));
 sky130_fd_sc_hd__dfxtp_1 _29469_ (.CLK(clknet_leaf_198_clk),
    .D(_00112_),
    .Q(\genblk1.pcpi_mul.rd[8] ));
 sky130_fd_sc_hd__dfxtp_1 _29470_ (.CLK(clknet_leaf_202_clk),
    .D(_00113_),
    .Q(\genblk1.pcpi_mul.rd[9] ));
 sky130_fd_sc_hd__dfxtp_1 _29471_ (.CLK(clknet_leaf_201_clk),
    .D(_00056_),
    .Q(\genblk1.pcpi_mul.rd[10] ));
 sky130_fd_sc_hd__dfxtp_1 _29472_ (.CLK(clknet_leaf_202_clk),
    .D(_00057_),
    .Q(\genblk1.pcpi_mul.rd[11] ));
 sky130_fd_sc_hd__dfxtp_1 _29473_ (.CLK(clknet_leaf_202_clk),
    .D(_00058_),
    .Q(\genblk1.pcpi_mul.rd[12] ));
 sky130_fd_sc_hd__dfxtp_1 _29474_ (.CLK(clknet_leaf_202_clk),
    .D(_00059_),
    .Q(\genblk1.pcpi_mul.rd[13] ));
 sky130_fd_sc_hd__dfxtp_1 _29475_ (.CLK(clknet_leaf_203_clk),
    .D(_00060_),
    .Q(\genblk1.pcpi_mul.rd[14] ));
 sky130_fd_sc_hd__dfxtp_1 _29476_ (.CLK(clknet_leaf_202_clk),
    .D(_00061_),
    .Q(\genblk1.pcpi_mul.rd[15] ));
 sky130_fd_sc_hd__dfxtp_1 _29477_ (.CLK(clknet_leaf_211_clk),
    .D(_00062_),
    .Q(\genblk1.pcpi_mul.rd[16] ));
 sky130_fd_sc_hd__dfxtp_1 _29478_ (.CLK(clknet_leaf_211_clk),
    .D(_00063_),
    .Q(\genblk1.pcpi_mul.rd[17] ));
 sky130_fd_sc_hd__dfxtp_1 _29479_ (.CLK(clknet_leaf_210_clk),
    .D(_00064_),
    .Q(\genblk1.pcpi_mul.rd[18] ));
 sky130_fd_sc_hd__dfxtp_1 _29480_ (.CLK(clknet_leaf_210_clk),
    .D(_00065_),
    .Q(\genblk1.pcpi_mul.rd[19] ));
 sky130_fd_sc_hd__dfxtp_1 _29481_ (.CLK(clknet_leaf_211_clk),
    .D(_00066_),
    .Q(\genblk1.pcpi_mul.rd[20] ));
 sky130_fd_sc_hd__dfxtp_1 _29482_ (.CLK(clknet_leaf_209_clk),
    .D(_00067_),
    .Q(\genblk1.pcpi_mul.rd[21] ));
 sky130_fd_sc_hd__dfxtp_1 _29483_ (.CLK(clknet_leaf_209_clk),
    .D(_00068_),
    .Q(\genblk1.pcpi_mul.rd[22] ));
 sky130_fd_sc_hd__dfxtp_1 _29484_ (.CLK(clknet_leaf_212_clk),
    .D(_00069_),
    .Q(\genblk1.pcpi_mul.rd[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29485_ (.CLK(clknet_5_0__leaf_clk),
    .D(_00070_),
    .Q(\genblk1.pcpi_mul.rd[24] ));
 sky130_fd_sc_hd__dfxtp_2 _29486_ (.CLK(clknet_leaf_3_clk),
    .D(_00071_),
    .Q(\genblk1.pcpi_mul.rd[25] ));
 sky130_fd_sc_hd__dfxtp_1 _29487_ (.CLK(clknet_leaf_4_clk),
    .D(_00072_),
    .Q(\genblk1.pcpi_mul.rd[26] ));
 sky130_fd_sc_hd__dfxtp_1 _29488_ (.CLK(clknet_leaf_3_clk),
    .D(_00073_),
    .Q(\genblk1.pcpi_mul.rd[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29489_ (.CLK(clknet_leaf_4_clk),
    .D(_00074_),
    .Q(\genblk1.pcpi_mul.rd[28] ));
 sky130_fd_sc_hd__dfxtp_2 _29490_ (.CLK(clknet_leaf_4_clk),
    .D(_00075_),
    .Q(\genblk1.pcpi_mul.rd[29] ));
 sky130_fd_sc_hd__dfxtp_2 _29491_ (.CLK(clknet_leaf_4_clk),
    .D(_00076_),
    .Q(\genblk1.pcpi_mul.rd[30] ));
 sky130_fd_sc_hd__dfxtp_2 _29492_ (.CLK(clknet_leaf_4_clk),
    .D(_00077_),
    .Q(\genblk1.pcpi_mul.rd[31] ));
 sky130_fd_sc_hd__dfxtp_1 _29493_ (.CLK(clknet_leaf_212_clk),
    .D(_00078_),
    .Q(\genblk1.pcpi_mul.rd[32] ));
 sky130_fd_sc_hd__dfxtp_1 _29494_ (.CLK(clknet_leaf_211_clk),
    .D(_00079_),
    .Q(\genblk1.pcpi_mul.rd[33] ));
 sky130_fd_sc_hd__dfxtp_1 _29495_ (.CLK(clknet_leaf_211_clk),
    .D(_00080_),
    .Q(\genblk1.pcpi_mul.rd[34] ));
 sky130_fd_sc_hd__dfxtp_1 _29496_ (.CLK(clknet_leaf_211_clk),
    .D(_00081_),
    .Q(\genblk1.pcpi_mul.rd[35] ));
 sky130_fd_sc_hd__dfxtp_1 _29497_ (.CLK(clknet_leaf_202_clk),
    .D(_00082_),
    .Q(\genblk1.pcpi_mul.rd[36] ));
 sky130_fd_sc_hd__dfxtp_1 _29498_ (.CLK(clknet_leaf_200_clk),
    .D(_00083_),
    .Q(\genblk1.pcpi_mul.rd[37] ));
 sky130_fd_sc_hd__dfxtp_1 _29499_ (.CLK(clknet_leaf_201_clk),
    .D(_00084_),
    .Q(\genblk1.pcpi_mul.rd[38] ));
 sky130_fd_sc_hd__dfxtp_1 _29500_ (.CLK(clknet_leaf_200_clk),
    .D(_00085_),
    .Q(\genblk1.pcpi_mul.rd[39] ));
 sky130_fd_sc_hd__dfxtp_1 _29501_ (.CLK(clknet_leaf_200_clk),
    .D(_00086_),
    .Q(\genblk1.pcpi_mul.rd[40] ));
 sky130_fd_sc_hd__dfxtp_1 _29502_ (.CLK(clknet_leaf_200_clk),
    .D(_00087_),
    .Q(\genblk1.pcpi_mul.rd[41] ));
 sky130_fd_sc_hd__dfxtp_1 _29503_ (.CLK(clknet_leaf_201_clk),
    .D(_00088_),
    .Q(\genblk1.pcpi_mul.rd[42] ));
 sky130_fd_sc_hd__dfxtp_1 _29504_ (.CLK(clknet_leaf_201_clk),
    .D(_00089_),
    .Q(\genblk1.pcpi_mul.rd[43] ));
 sky130_fd_sc_hd__dfxtp_1 _29505_ (.CLK(clknet_leaf_200_clk),
    .D(_00090_),
    .Q(\genblk1.pcpi_mul.rd[44] ));
 sky130_fd_sc_hd__dfxtp_1 _29506_ (.CLK(clknet_leaf_200_clk),
    .D(_00091_),
    .Q(\genblk1.pcpi_mul.rd[45] ));
 sky130_fd_sc_hd__dfxtp_1 _29507_ (.CLK(clknet_leaf_200_clk),
    .D(_00092_),
    .Q(\genblk1.pcpi_mul.rd[46] ));
 sky130_fd_sc_hd__dfxtp_1 _29508_ (.CLK(clknet_leaf_201_clk),
    .D(_00093_),
    .Q(\genblk1.pcpi_mul.rd[47] ));
 sky130_fd_sc_hd__dfxtp_1 _29509_ (.CLK(clknet_leaf_202_clk),
    .D(_00094_),
    .Q(\genblk1.pcpi_mul.rd[48] ));
 sky130_fd_sc_hd__dfxtp_1 _29510_ (.CLK(clknet_leaf_201_clk),
    .D(_00095_),
    .Q(\genblk1.pcpi_mul.rd[49] ));
 sky130_fd_sc_hd__dfxtp_1 _29511_ (.CLK(clknet_leaf_201_clk),
    .D(_00096_),
    .Q(\genblk1.pcpi_mul.rd[50] ));
 sky130_fd_sc_hd__dfxtp_1 _29512_ (.CLK(clknet_leaf_201_clk),
    .D(_00097_),
    .Q(\genblk1.pcpi_mul.rd[51] ));
 sky130_fd_sc_hd__dfxtp_1 _29513_ (.CLK(clknet_leaf_201_clk),
    .D(_00098_),
    .Q(\genblk1.pcpi_mul.rd[52] ));
 sky130_fd_sc_hd__dfxtp_1 _29514_ (.CLK(clknet_leaf_201_clk),
    .D(_00099_),
    .Q(\genblk1.pcpi_mul.rd[53] ));
 sky130_fd_sc_hd__dfxtp_1 _29515_ (.CLK(clknet_leaf_201_clk),
    .D(_00100_),
    .Q(\genblk1.pcpi_mul.rd[54] ));
 sky130_fd_sc_hd__dfxtp_1 _29516_ (.CLK(clknet_leaf_201_clk),
    .D(_00101_),
    .Q(\genblk1.pcpi_mul.rd[55] ));
 sky130_fd_sc_hd__dfxtp_1 _29517_ (.CLK(clknet_leaf_202_clk),
    .D(_00102_),
    .Q(\genblk1.pcpi_mul.rd[56] ));
 sky130_fd_sc_hd__dfxtp_2 _29518_ (.CLK(clknet_leaf_195_clk),
    .D(_00103_),
    .Q(\genblk1.pcpi_mul.rd[57] ));
 sky130_fd_sc_hd__dfxtp_2 _29519_ (.CLK(clknet_leaf_195_clk),
    .D(_00104_),
    .Q(\genblk1.pcpi_mul.rd[58] ));
 sky130_fd_sc_hd__dfxtp_2 _29520_ (.CLK(clknet_leaf_195_clk),
    .D(_00105_),
    .Q(\genblk1.pcpi_mul.rd[59] ));
 sky130_fd_sc_hd__dfxtp_2 _29521_ (.CLK(clknet_leaf_195_clk),
    .D(_00106_),
    .Q(\genblk1.pcpi_mul.rd[60] ));
 sky130_fd_sc_hd__dfxtp_2 _29522_ (.CLK(clknet_leaf_195_clk),
    .D(_00107_),
    .Q(\genblk1.pcpi_mul.rd[61] ));
 sky130_fd_sc_hd__dfxtp_2 _29523_ (.CLK(clknet_leaf_194_clk),
    .D(_00108_),
    .Q(\genblk1.pcpi_mul.rd[62] ));
 sky130_fd_sc_hd__dfxtp_2 _29524_ (.CLK(clknet_leaf_194_clk),
    .D(_00109_),
    .Q(\genblk1.pcpi_mul.rd[63] ));
 sky130_fd_sc_hd__dfxtp_1 _29525_ (.CLK(clknet_leaf_186_clk),
    .D(_00178_),
    .Q(\cpuregs[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29526_ (.CLK(clknet_leaf_181_clk),
    .D(_00179_),
    .Q(\cpuregs[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29527_ (.CLK(clknet_leaf_180_clk),
    .D(_00180_),
    .Q(\cpuregs[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29528_ (.CLK(clknet_leaf_180_clk),
    .D(_00181_),
    .Q(\cpuregs[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29529_ (.CLK(clknet_leaf_179_clk),
    .D(_00182_),
    .Q(\cpuregs[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29530_ (.CLK(clknet_leaf_185_clk),
    .D(_00183_),
    .Q(\cpuregs[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29531_ (.CLK(clknet_leaf_183_clk),
    .D(_00184_),
    .Q(\cpuregs[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29532_ (.CLK(clknet_leaf_191_clk),
    .D(_00185_),
    .Q(\cpuregs[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29533_ (.CLK(clknet_leaf_191_clk),
    .D(_00186_),
    .Q(\cpuregs[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29534_ (.CLK(clknet_leaf_188_clk),
    .D(_00187_),
    .Q(\cpuregs[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29535_ (.CLK(clknet_leaf_189_clk),
    .D(_00188_),
    .Q(\cpuregs[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29536_ (.CLK(clknet_leaf_183_clk),
    .D(_00189_),
    .Q(\cpuregs[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29537_ (.CLK(clknet_leaf_124_clk),
    .D(_00190_),
    .Q(\cpuregs[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29538_ (.CLK(clknet_leaf_100_clk),
    .D(_00191_),
    .Q(\cpuregs[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29539_ (.CLK(clknet_leaf_99_clk),
    .D(_00192_),
    .Q(\cpuregs[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29540_ (.CLK(clknet_leaf_140_clk),
    .D(_00193_),
    .Q(\cpuregs[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29541_ (.CLK(clknet_leaf_124_clk),
    .D(_00194_),
    .Q(\cpuregs[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29542_ (.CLK(clknet_leaf_101_clk),
    .D(_00195_),
    .Q(\cpuregs[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29543_ (.CLK(clknet_leaf_154_clk),
    .D(_00196_),
    .Q(\cpuregs[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29544_ (.CLK(clknet_leaf_157_clk),
    .D(_00197_),
    .Q(\cpuregs[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29545_ (.CLK(clknet_leaf_155_clk),
    .D(_00198_),
    .Q(\cpuregs[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29546_ (.CLK(clknet_leaf_160_clk),
    .D(_00199_),
    .Q(\cpuregs[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29547_ (.CLK(clknet_leaf_154_clk),
    .D(_00200_),
    .Q(\cpuregs[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29548_ (.CLK(clknet_leaf_155_clk),
    .D(_00201_),
    .Q(\cpuregs[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29549_ (.CLK(clknet_leaf_129_clk),
    .D(_00202_),
    .Q(\cpuregs[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29550_ (.CLK(clknet_leaf_130_clk),
    .D(_00203_),
    .Q(\cpuregs[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29551_ (.CLK(clknet_leaf_126_clk),
    .D(_00204_),
    .Q(\cpuregs[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29552_ (.CLK(clknet_leaf_126_clk),
    .D(_00205_),
    .Q(\cpuregs[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29553_ (.CLK(clknet_leaf_125_clk),
    .D(_00206_),
    .Q(\cpuregs[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29554_ (.CLK(clknet_leaf_127_clk),
    .D(_00207_),
    .Q(\cpuregs[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29555_ (.CLK(clknet_leaf_133_clk),
    .D(_00208_),
    .Q(\cpuregs[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29556_ (.CLK(clknet_leaf_145_clk),
    .D(_00209_),
    .Q(\cpuregs[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29557_ (.CLK(clknet_leaf_187_clk),
    .D(_00210_),
    .Q(\cpuregs[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29558_ (.CLK(clknet_leaf_181_clk),
    .D(_00211_),
    .Q(\cpuregs[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29559_ (.CLK(clknet_leaf_180_clk),
    .D(_00212_),
    .Q(\cpuregs[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29560_ (.CLK(clknet_leaf_179_clk),
    .D(_00213_),
    .Q(\cpuregs[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29561_ (.CLK(clknet_leaf_179_clk),
    .D(_00214_),
    .Q(\cpuregs[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29562_ (.CLK(clknet_leaf_185_clk),
    .D(_00215_),
    .Q(\cpuregs[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29563_ (.CLK(clknet_leaf_184_clk),
    .D(_00216_),
    .Q(\cpuregs[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29564_ (.CLK(clknet_leaf_194_clk),
    .D(_00217_),
    .Q(\cpuregs[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29565_ (.CLK(clknet_leaf_191_clk),
    .D(_00218_),
    .Q(\cpuregs[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29566_ (.CLK(clknet_leaf_188_clk),
    .D(_00219_),
    .Q(\cpuregs[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29567_ (.CLK(clknet_leaf_190_clk),
    .D(_00220_),
    .Q(\cpuregs[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29568_ (.CLK(clknet_leaf_183_clk),
    .D(_00221_),
    .Q(\cpuregs[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29569_ (.CLK(clknet_leaf_139_clk),
    .D(_00222_),
    .Q(\cpuregs[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29570_ (.CLK(clknet_leaf_100_clk),
    .D(_00223_),
    .Q(\cpuregs[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29571_ (.CLK(clknet_leaf_100_clk),
    .D(_00224_),
    .Q(\cpuregs[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29572_ (.CLK(clknet_leaf_139_clk),
    .D(_00225_),
    .Q(\cpuregs[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29573_ (.CLK(clknet_leaf_139_clk),
    .D(_00226_),
    .Q(\cpuregs[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29574_ (.CLK(clknet_leaf_122_clk),
    .D(_00227_),
    .Q(\cpuregs[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29575_ (.CLK(clknet_leaf_154_clk),
    .D(_00228_),
    .Q(\cpuregs[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29576_ (.CLK(clknet_leaf_155_clk),
    .D(_00229_),
    .Q(\cpuregs[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29577_ (.CLK(clknet_leaf_149_clk),
    .D(_00230_),
    .Q(\cpuregs[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29578_ (.CLK(clknet_leaf_150_clk),
    .D(_00231_),
    .Q(\cpuregs[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29579_ (.CLK(clknet_leaf_151_clk),
    .D(_00232_),
    .Q(\cpuregs[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29580_ (.CLK(clknet_leaf_155_clk),
    .D(_00233_),
    .Q(\cpuregs[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29581_ (.CLK(clknet_leaf_129_clk),
    .D(_00234_),
    .Q(\cpuregs[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29582_ (.CLK(clknet_leaf_129_clk),
    .D(_00235_),
    .Q(\cpuregs[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29583_ (.CLK(clknet_leaf_126_clk),
    .D(_00236_),
    .Q(\cpuregs[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29584_ (.CLK(clknet_leaf_127_clk),
    .D(_00237_),
    .Q(\cpuregs[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29585_ (.CLK(clknet_leaf_129_clk),
    .D(_00238_),
    .Q(\cpuregs[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29586_ (.CLK(clknet_leaf_127_clk),
    .D(_00239_),
    .Q(\cpuregs[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29587_ (.CLK(clknet_leaf_133_clk),
    .D(_00240_),
    .Q(\cpuregs[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29588_ (.CLK(clknet_leaf_145_clk),
    .D(_00241_),
    .Q(\cpuregs[6][31] ));
 sky130_fd_sc_hd__dfxtp_2 _29589_ (.CLK(clknet_leaf_17_clk),
    .D(_00242_),
    .Q(\genblk1.pcpi_mul.rs2[32] ));
 sky130_fd_sc_hd__dfxtp_4 _29590_ (.CLK(clknet_leaf_17_clk),
    .D(_00243_),
    .Q(\genblk1.pcpi_mul.rs1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _29591_ (.CLK(clknet_leaf_158_clk),
    .D(_00244_),
    .Q(\cpuregs[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29592_ (.CLK(clknet_leaf_179_clk),
    .D(_00245_),
    .Q(\cpuregs[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29593_ (.CLK(clknet_leaf_180_clk),
    .D(_00246_),
    .Q(\cpuregs[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29594_ (.CLK(clknet_leaf_185_clk),
    .D(_00247_),
    .Q(\cpuregs[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29595_ (.CLK(clknet_leaf_179_clk),
    .D(_00248_),
    .Q(\cpuregs[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29596_ (.CLK(clknet_leaf_158_clk),
    .D(_00249_),
    .Q(\cpuregs[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29597_ (.CLK(clknet_leaf_184_clk),
    .D(_00250_),
    .Q(\cpuregs[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29598_ (.CLK(clknet_leaf_194_clk),
    .D(_00251_),
    .Q(\cpuregs[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29599_ (.CLK(clknet_leaf_191_clk),
    .D(_00252_),
    .Q(\cpuregs[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29600_ (.CLK(clknet_leaf_191_clk),
    .D(_00253_),
    .Q(\cpuregs[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29601_ (.CLK(clknet_leaf_194_clk),
    .D(_00254_),
    .Q(\cpuregs[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29602_ (.CLK(clknet_leaf_183_clk),
    .D(_00255_),
    .Q(\cpuregs[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29603_ (.CLK(clknet_leaf_139_clk),
    .D(_00256_),
    .Q(\cpuregs[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29604_ (.CLK(clknet_leaf_122_clk),
    .D(_00257_),
    .Q(\cpuregs[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29605_ (.CLK(clknet_leaf_100_clk),
    .D(_00258_),
    .Q(\cpuregs[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29606_ (.CLK(clknet_leaf_139_clk),
    .D(_00259_),
    .Q(\cpuregs[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29607_ (.CLK(clknet_leaf_139_clk),
    .D(_00260_),
    .Q(\cpuregs[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29608_ (.CLK(clknet_leaf_122_clk),
    .D(_00261_),
    .Q(\cpuregs[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29609_ (.CLK(clknet_leaf_153_clk),
    .D(_00262_),
    .Q(\cpuregs[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29610_ (.CLK(clknet_leaf_154_clk),
    .D(_00263_),
    .Q(\cpuregs[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29611_ (.CLK(clknet_leaf_154_clk),
    .D(_00264_),
    .Q(\cpuregs[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29612_ (.CLK(clknet_leaf_151_clk),
    .D(_00265_),
    .Q(\cpuregs[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29613_ (.CLK(clknet_leaf_151_clk),
    .D(_00266_),
    .Q(\cpuregs[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29614_ (.CLK(clknet_leaf_154_clk),
    .D(_00267_),
    .Q(\cpuregs[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29615_ (.CLK(clknet_leaf_129_clk),
    .D(_00268_),
    .Q(\cpuregs[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29616_ (.CLK(clknet_leaf_130_clk),
    .D(_00269_),
    .Q(\cpuregs[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29617_ (.CLK(clknet_leaf_127_clk),
    .D(_00270_),
    .Q(\cpuregs[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29618_ (.CLK(clknet_leaf_127_clk),
    .D(_00271_),
    .Q(\cpuregs[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29619_ (.CLK(clknet_leaf_129_clk),
    .D(_00272_),
    .Q(\cpuregs[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29620_ (.CLK(clknet_leaf_127_clk),
    .D(_00273_),
    .Q(\cpuregs[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29621_ (.CLK(clknet_leaf_132_clk),
    .D(_00274_),
    .Q(\cpuregs[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29622_ (.CLK(clknet_leaf_146_clk),
    .D(_00275_),
    .Q(\cpuregs[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29623_ (.CLK(clknet_leaf_157_clk),
    .D(_00276_),
    .Q(\cpuregs[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29624_ (.CLK(clknet_leaf_177_clk),
    .D(_00277_),
    .Q(\cpuregs[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29625_ (.CLK(clknet_leaf_177_clk),
    .D(_00278_),
    .Q(\cpuregs[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29626_ (.CLK(clknet_leaf_186_clk),
    .D(_00279_),
    .Q(\cpuregs[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29627_ (.CLK(clknet_leaf_178_clk),
    .D(_00280_),
    .Q(\cpuregs[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29628_ (.CLK(clknet_leaf_169_clk),
    .D(_00281_),
    .Q(\cpuregs[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29629_ (.CLK(clknet_leaf_186_clk),
    .D(_00282_),
    .Q(\cpuregs[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29630_ (.CLK(clknet_leaf_190_clk),
    .D(_00283_),
    .Q(\cpuregs[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29631_ (.CLK(clknet_leaf_156_clk),
    .D(_00284_),
    .Q(\cpuregs[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29632_ (.CLK(clknet_leaf_154_clk),
    .D(_00285_),
    .Q(\cpuregs[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29633_ (.CLK(clknet_leaf_189_clk),
    .D(_00286_),
    .Q(\cpuregs[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29634_ (.CLK(clknet_leaf_189_clk),
    .D(_00287_),
    .Q(\cpuregs[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29635_ (.CLK(clknet_leaf_139_clk),
    .D(_00288_),
    .Q(\cpuregs[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29636_ (.CLK(clknet_leaf_140_clk),
    .D(_00289_),
    .Q(\cpuregs[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29637_ (.CLK(clknet_leaf_100_clk),
    .D(_00290_),
    .Q(\cpuregs[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29638_ (.CLK(clknet_leaf_141_clk),
    .D(_00291_),
    .Q(\cpuregs[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29639_ (.CLK(clknet_leaf_137_clk),
    .D(_00292_),
    .Q(\cpuregs[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29640_ (.CLK(clknet_leaf_122_clk),
    .D(_00293_),
    .Q(\cpuregs[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29641_ (.CLK(clknet_leaf_161_clk),
    .D(_00294_),
    .Q(\cpuregs[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29642_ (.CLK(clknet_leaf_149_clk),
    .D(_00295_),
    .Q(\cpuregs[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29643_ (.CLK(clknet_leaf_149_clk),
    .D(_00296_),
    .Q(\cpuregs[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29644_ (.CLK(clknet_leaf_148_clk),
    .D(_00297_),
    .Q(\cpuregs[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29645_ (.CLK(clknet_leaf_148_clk),
    .D(_00298_),
    .Q(\cpuregs[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29646_ (.CLK(clknet_leaf_161_clk),
    .D(_00299_),
    .Q(\cpuregs[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29647_ (.CLK(clknet_leaf_130_clk),
    .D(_00300_),
    .Q(\cpuregs[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29648_ (.CLK(clknet_leaf_132_clk),
    .D(_00301_),
    .Q(\cpuregs[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29649_ (.CLK(clknet_leaf_121_clk),
    .D(_00302_),
    .Q(\cpuregs[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29650_ (.CLK(clknet_leaf_118_clk),
    .D(_00303_),
    .Q(\cpuregs[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29651_ (.CLK(clknet_leaf_126_clk),
    .D(_00304_),
    .Q(\cpuregs[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29652_ (.CLK(clknet_leaf_118_clk),
    .D(_00305_),
    .Q(\cpuregs[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29653_ (.CLK(clknet_leaf_138_clk),
    .D(_00306_),
    .Q(\cpuregs[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29654_ (.CLK(clknet_leaf_142_clk),
    .D(_00307_),
    .Q(\cpuregs[8][31] ));
 sky130_fd_sc_hd__dfxtp_2 _29655_ (.CLK(clknet_leaf_30_clk),
    .D(_00308_),
    .Q(\decoded_imm_uj[4] ));
 sky130_fd_sc_hd__dfxtp_2 _29656_ (.CLK(clknet_leaf_30_clk),
    .D(_00309_),
    .Q(\decoded_imm_uj[5] ));
 sky130_fd_sc_hd__dfxtp_1 _29657_ (.CLK(clknet_leaf_29_clk),
    .D(_00310_),
    .Q(\decoded_imm_uj[6] ));
 sky130_fd_sc_hd__dfxtp_1 _29658_ (.CLK(clknet_leaf_30_clk),
    .D(_00311_),
    .Q(\decoded_imm_uj[7] ));
 sky130_fd_sc_hd__dfxtp_1 _29659_ (.CLK(clknet_leaf_29_clk),
    .D(_00312_),
    .Q(\decoded_imm_uj[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29660_ (.CLK(clknet_leaf_28_clk),
    .D(_00313_),
    .Q(\decoded_imm_uj[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29661_ (.CLK(clknet_leaf_27_clk),
    .D(_00314_),
    .Q(\decoded_imm_uj[10] ));
 sky130_fd_sc_hd__dfxtp_1 _29662_ (.CLK(clknet_leaf_26_clk),
    .D(_00315_),
    .Q(\decoded_imm_uj[12] ));
 sky130_fd_sc_hd__dfxtp_1 _29663_ (.CLK(clknet_leaf_26_clk),
    .D(_00316_),
    .Q(\decoded_imm_uj[13] ));
 sky130_fd_sc_hd__dfxtp_1 _29664_ (.CLK(clknet_leaf_26_clk),
    .D(_00317_),
    .Q(\decoded_imm_uj[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29665_ (.CLK(clknet_leaf_95_clk),
    .D(_00318_),
    .Q(\decoded_imm_uj[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29666_ (.CLK(clknet_leaf_95_clk),
    .D(_00319_),
    .Q(\decoded_imm_uj[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29667_ (.CLK(clknet_leaf_95_clk),
    .D(_00320_),
    .Q(\decoded_imm_uj[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29668_ (.CLK(clknet_leaf_95_clk),
    .D(_00321_),
    .Q(\decoded_imm_uj[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29669_ (.CLK(clknet_leaf_24_clk),
    .D(_00322_),
    .Q(\decoded_imm_uj[19] ));
 sky130_fd_sc_hd__dfxtp_2 _29670_ (.CLK(clknet_leaf_176_clk),
    .D(_00323_),
    .Q(\decoded_imm_uj[20] ));
 sky130_fd_sc_hd__dfxtp_1 _29671_ (.CLK(clknet_leaf_160_clk),
    .D(_00324_),
    .Q(\cpuregs[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29672_ (.CLK(clknet_leaf_181_clk),
    .D(_00325_),
    .Q(\cpuregs[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29673_ (.CLK(clknet_leaf_172_clk),
    .D(_00326_),
    .Q(\cpuregs[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29674_ (.CLK(clknet_leaf_160_clk),
    .D(_00327_),
    .Q(\cpuregs[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29675_ (.CLK(clknet_leaf_170_clk),
    .D(_00328_),
    .Q(\cpuregs[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29676_ (.CLK(clknet_leaf_169_clk),
    .D(_00329_),
    .Q(\cpuregs[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29677_ (.CLK(clknet_leaf_185_clk),
    .D(_00330_),
    .Q(\cpuregs[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29678_ (.CLK(clknet_leaf_193_clk),
    .D(_00331_),
    .Q(\cpuregs[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29679_ (.CLK(clknet_leaf_192_clk),
    .D(_00332_),
    .Q(\cpuregs[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29680_ (.CLK(clknet_leaf_152_clk),
    .D(_00333_),
    .Q(\cpuregs[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29681_ (.CLK(clknet_leaf_183_clk),
    .D(_00334_),
    .Q(\cpuregs[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29682_ (.CLK(clknet_leaf_156_clk),
    .D(_00335_),
    .Q(\cpuregs[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29683_ (.CLK(clknet_leaf_139_clk),
    .D(_00336_),
    .Q(\cpuregs[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29684_ (.CLK(clknet_leaf_122_clk),
    .D(_00337_),
    .Q(\cpuregs[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29685_ (.CLK(clknet_leaf_165_clk),
    .D(_00338_),
    .Q(\cpuregs[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29686_ (.CLK(clknet_leaf_164_clk),
    .D(_00339_),
    .Q(\cpuregs[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29687_ (.CLK(clknet_leaf_134_clk),
    .D(_00340_),
    .Q(\cpuregs[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29688_ (.CLK(clknet_leaf_121_clk),
    .D(_00341_),
    .Q(\cpuregs[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29689_ (.CLK(clknet_leaf_142_clk),
    .D(_00342_),
    .Q(\cpuregs[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29690_ (.CLK(clknet_leaf_163_clk),
    .D(_00343_),
    .Q(\cpuregs[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29691_ (.CLK(clknet_leaf_162_clk),
    .D(_00344_),
    .Q(\cpuregs[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29692_ (.CLK(clknet_leaf_162_clk),
    .D(_00345_),
    .Q(\cpuregs[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29693_ (.CLK(clknet_leaf_142_clk),
    .D(_00346_),
    .Q(\cpuregs[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29694_ (.CLK(clknet_leaf_160_clk),
    .D(_00347_),
    .Q(\cpuregs[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29695_ (.CLK(clknet_leaf_123_clk),
    .D(_00348_),
    .Q(\cpuregs[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29696_ (.CLK(clknet_leaf_138_clk),
    .D(_00349_),
    .Q(\cpuregs[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29697_ (.CLK(clknet_leaf_117_clk),
    .D(_00350_),
    .Q(\cpuregs[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29698_ (.CLK(clknet_leaf_119_clk),
    .D(_00351_),
    .Q(\cpuregs[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29699_ (.CLK(clknet_leaf_125_clk),
    .D(_00352_),
    .Q(\cpuregs[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29700_ (.CLK(clknet_leaf_116_clk),
    .D(_00353_),
    .Q(\cpuregs[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29701_ (.CLK(clknet_leaf_134_clk),
    .D(_00354_),
    .Q(\cpuregs[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29702_ (.CLK(clknet_leaf_142_clk),
    .D(_00355_),
    .Q(\cpuregs[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29703_ (.CLK(clknet_leaf_157_clk),
    .D(_00356_),
    .Q(\cpuregs[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29704_ (.CLK(clknet_leaf_181_clk),
    .D(_00357_),
    .Q(\cpuregs[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29705_ (.CLK(clknet_leaf_181_clk),
    .D(_00358_),
    .Q(\cpuregs[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29706_ (.CLK(clknet_leaf_186_clk),
    .D(_00359_),
    .Q(\cpuregs[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29707_ (.CLK(clknet_leaf_179_clk),
    .D(_00360_),
    .Q(\cpuregs[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29708_ (.CLK(clknet_leaf_170_clk),
    .D(_00361_),
    .Q(\cpuregs[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29709_ (.CLK(clknet_leaf_184_clk),
    .D(_00362_),
    .Q(\cpuregs[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29710_ (.CLK(clknet_leaf_194_clk),
    .D(_00363_),
    .Q(\cpuregs[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29711_ (.CLK(clknet_leaf_191_clk),
    .D(_00364_),
    .Q(\cpuregs[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29712_ (.CLK(clknet_leaf_188_clk),
    .D(_00365_),
    .Q(\cpuregs[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29713_ (.CLK(clknet_leaf_190_clk),
    .D(_00366_),
    .Q(\cpuregs[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29714_ (.CLK(clknet_leaf_183_clk),
    .D(_00367_),
    .Q(\cpuregs[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29715_ (.CLK(clknet_leaf_139_clk),
    .D(_00368_),
    .Q(\cpuregs[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29716_ (.CLK(clknet_leaf_140_clk),
    .D(_00369_),
    .Q(\cpuregs[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29717_ (.CLK(clknet_leaf_123_clk),
    .D(_00370_),
    .Q(\cpuregs[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29718_ (.CLK(clknet_leaf_139_clk),
    .D(_00371_),
    .Q(\cpuregs[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29719_ (.CLK(clknet_leaf_139_clk),
    .D(_00372_),
    .Q(\cpuregs[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29720_ (.CLK(clknet_leaf_122_clk),
    .D(_00373_),
    .Q(\cpuregs[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29721_ (.CLK(clknet_leaf_150_clk),
    .D(_00374_),
    .Q(\cpuregs[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29722_ (.CLK(clknet_leaf_149_clk),
    .D(_00375_),
    .Q(\cpuregs[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29723_ (.CLK(clknet_leaf_149_clk),
    .D(_00376_),
    .Q(\cpuregs[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29724_ (.CLK(clknet_leaf_150_clk),
    .D(_00377_),
    .Q(\cpuregs[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29725_ (.CLK(clknet_leaf_148_clk),
    .D(_00378_),
    .Q(\cpuregs[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29726_ (.CLK(clknet_leaf_161_clk),
    .D(_00379_),
    .Q(\cpuregs[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29727_ (.CLK(clknet_leaf_130_clk),
    .D(_00380_),
    .Q(\cpuregs[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29728_ (.CLK(clknet_leaf_130_clk),
    .D(_00381_),
    .Q(\cpuregs[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29729_ (.CLK(clknet_leaf_127_clk),
    .D(_00382_),
    .Q(\cpuregs[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29730_ (.CLK(clknet_leaf_118_clk),
    .D(_00383_),
    .Q(\cpuregs[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29731_ (.CLK(clknet_leaf_127_clk),
    .D(_00384_),
    .Q(\cpuregs[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29732_ (.CLK(clknet_leaf_118_clk),
    .D(_00385_),
    .Q(\cpuregs[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29733_ (.CLK(clknet_leaf_133_clk),
    .D(_00386_),
    .Q(\cpuregs[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29734_ (.CLK(clknet_leaf_145_clk),
    .D(_00387_),
    .Q(\cpuregs[10][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29735_ (.CLK(clknet_leaf_212_clk),
    .D(\genblk1.pcpi_mul.instr_any_mulh ),
    .Q(\genblk1.pcpi_mul.shift_out ));
 sky130_fd_sc_hd__dfxtp_1 _29736_ (.CLK(clknet_leaf_157_clk),
    .D(_00388_),
    .Q(\cpuregs[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29737_ (.CLK(clknet_leaf_181_clk),
    .D(_00389_),
    .Q(\cpuregs[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29738_ (.CLK(clknet_leaf_177_clk),
    .D(_00390_),
    .Q(\cpuregs[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29739_ (.CLK(clknet_leaf_185_clk),
    .D(_00391_),
    .Q(\cpuregs[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29740_ (.CLK(clknet_leaf_178_clk),
    .D(_00392_),
    .Q(\cpuregs[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29741_ (.CLK(clknet_leaf_169_clk),
    .D(_00393_),
    .Q(\cpuregs[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29742_ (.CLK(clknet_leaf_183_clk),
    .D(_00394_),
    .Q(\cpuregs[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29743_ (.CLK(clknet_leaf_193_clk),
    .D(_00395_),
    .Q(\cpuregs[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29744_ (.CLK(clknet_leaf_191_clk),
    .D(_00396_),
    .Q(\cpuregs[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29745_ (.CLK(clknet_leaf_191_clk),
    .D(_00397_),
    .Q(\cpuregs[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29746_ (.CLK(clknet_leaf_194_clk),
    .D(_00398_),
    .Q(\cpuregs[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29747_ (.CLK(clknet_leaf_183_clk),
    .D(_00399_),
    .Q(\cpuregs[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29748_ (.CLK(clknet_leaf_137_clk),
    .D(_00400_),
    .Q(\cpuregs[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29749_ (.CLK(clknet_leaf_140_clk),
    .D(_00401_),
    .Q(\cpuregs[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29750_ (.CLK(clknet_leaf_123_clk),
    .D(_00402_),
    .Q(\cpuregs[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29751_ (.CLK(clknet_leaf_137_clk),
    .D(_00403_),
    .Q(\cpuregs[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29752_ (.CLK(clknet_leaf_137_clk),
    .D(_00404_),
    .Q(\cpuregs[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29753_ (.CLK(clknet_leaf_123_clk),
    .D(_00405_),
    .Q(\cpuregs[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29754_ (.CLK(clknet_leaf_150_clk),
    .D(_00406_),
    .Q(\cpuregs[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29755_ (.CLK(clknet_leaf_151_clk),
    .D(_00407_),
    .Q(\cpuregs[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29756_ (.CLK(clknet_leaf_149_clk),
    .D(_00408_),
    .Q(\cpuregs[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29757_ (.CLK(clknet_leaf_151_clk),
    .D(_00409_),
    .Q(\cpuregs[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29758_ (.CLK(clknet_leaf_148_clk),
    .D(_00410_),
    .Q(\cpuregs[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29759_ (.CLK(clknet_leaf_150_clk),
    .D(_00411_),
    .Q(\cpuregs[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29760_ (.CLK(clknet_5_31__leaf_clk),
    .D(_00412_),
    .Q(\cpuregs[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29761_ (.CLK(clknet_leaf_130_clk),
    .D(_00413_),
    .Q(\cpuregs[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29762_ (.CLK(clknet_leaf_128_clk),
    .D(_00414_),
    .Q(\cpuregs[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29763_ (.CLK(clknet_leaf_117_clk),
    .D(_00415_),
    .Q(\cpuregs[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29764_ (.CLK(clknet_leaf_126_clk),
    .D(_00416_),
    .Q(\cpuregs[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29765_ (.CLK(clknet_leaf_117_clk),
    .D(_00417_),
    .Q(\cpuregs[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29766_ (.CLK(clknet_leaf_133_clk),
    .D(_00418_),
    .Q(\cpuregs[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29767_ (.CLK(clknet_leaf_145_clk),
    .D(_00419_),
    .Q(\cpuregs[11][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29768_ (.CLK(clknet_leaf_158_clk),
    .D(_00420_),
    .Q(\cpuregs[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29769_ (.CLK(clknet_leaf_177_clk),
    .D(_00421_),
    .Q(\cpuregs[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29770_ (.CLK(clknet_leaf_172_clk),
    .D(_00422_),
    .Q(\cpuregs[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29771_ (.CLK(clknet_leaf_158_clk),
    .D(_00423_),
    .Q(\cpuregs[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29772_ (.CLK(clknet_leaf_178_clk),
    .D(_00424_),
    .Q(\cpuregs[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29773_ (.CLK(clknet_leaf_169_clk),
    .D(_00425_),
    .Q(\cpuregs[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29774_ (.CLK(clknet_leaf_189_clk),
    .D(_00426_),
    .Q(\cpuregs[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29775_ (.CLK(clknet_leaf_193_clk),
    .D(_00427_),
    .Q(\cpuregs[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29776_ (.CLK(clknet_leaf_191_clk),
    .D(_00428_),
    .Q(\cpuregs[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29777_ (.CLK(clknet_leaf_153_clk),
    .D(_00429_),
    .Q(\cpuregs[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29778_ (.CLK(clknet_leaf_190_clk),
    .D(_00430_),
    .Q(\cpuregs[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29779_ (.CLK(clknet_leaf_156_clk),
    .D(_00431_),
    .Q(\cpuregs[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29780_ (.CLK(clknet_leaf_136_clk),
    .D(_00432_),
    .Q(\cpuregs[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29781_ (.CLK(clknet_leaf_141_clk),
    .D(_00433_),
    .Q(\cpuregs[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29782_ (.CLK(clknet_leaf_140_clk),
    .D(_00434_),
    .Q(\cpuregs[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29783_ (.CLK(clknet_leaf_136_clk),
    .D(_00435_),
    .Q(\cpuregs[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29784_ (.CLK(clknet_leaf_137_clk),
    .D(_00436_),
    .Q(\cpuregs[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29785_ (.CLK(clknet_leaf_123_clk),
    .D(_00437_),
    .Q(\cpuregs[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29786_ (.CLK(clknet_leaf_149_clk),
    .D(_00438_),
    .Q(\cpuregs[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29787_ (.CLK(clknet_leaf_147_clk),
    .D(_00439_),
    .Q(\cpuregs[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29788_ (.CLK(clknet_leaf_143_clk),
    .D(_00440_),
    .Q(\cpuregs[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29789_ (.CLK(clknet_leaf_147_clk),
    .D(_00441_),
    .Q(\cpuregs[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29790_ (.CLK(clknet_leaf_145_clk),
    .D(_00442_),
    .Q(\cpuregs[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29791_ (.CLK(clknet_leaf_161_clk),
    .D(_00443_),
    .Q(\cpuregs[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29792_ (.CLK(clknet_leaf_129_clk),
    .D(_00444_),
    .Q(\cpuregs[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29793_ (.CLK(clknet_leaf_130_clk),
    .D(_00445_),
    .Q(\cpuregs[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29794_ (.CLK(clknet_leaf_117_clk),
    .D(_00446_),
    .Q(\cpuregs[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29795_ (.CLK(clknet_leaf_118_clk),
    .D(_00447_),
    .Q(\cpuregs[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29796_ (.CLK(clknet_leaf_124_clk),
    .D(_00448_),
    .Q(\cpuregs[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29797_ (.CLK(clknet_leaf_119_clk),
    .D(_00449_),
    .Q(\cpuregs[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29798_ (.CLK(clknet_leaf_134_clk),
    .D(_00450_),
    .Q(\cpuregs[12][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29799_ (.CLK(clknet_leaf_145_clk),
    .D(_00451_),
    .Q(\cpuregs[12][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29800_ (.CLK(clknet_leaf_84_clk),
    .D(_00452_),
    .Q(net198));
 sky130_fd_sc_hd__dfxtp_1 _29801_ (.CLK(clknet_leaf_158_clk),
    .D(_00453_),
    .Q(\cpuregs[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29802_ (.CLK(clknet_leaf_177_clk),
    .D(_00454_),
    .Q(\cpuregs[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29803_ (.CLK(clknet_leaf_171_clk),
    .D(_00455_),
    .Q(\cpuregs[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29804_ (.CLK(clknet_leaf_156_clk),
    .D(_00456_),
    .Q(\cpuregs[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29805_ (.CLK(clknet_leaf_178_clk),
    .D(_00457_),
    .Q(\cpuregs[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29806_ (.CLK(clknet_leaf_169_clk),
    .D(_00458_),
    .Q(\cpuregs[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29807_ (.CLK(clknet_leaf_184_clk),
    .D(_00459_),
    .Q(\cpuregs[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29808_ (.CLK(clknet_leaf_193_clk),
    .D(_00460_),
    .Q(\cpuregs[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29809_ (.CLK(clknet_leaf_191_clk),
    .D(_00461_),
    .Q(\cpuregs[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29810_ (.CLK(clknet_leaf_153_clk),
    .D(_00462_),
    .Q(\cpuregs[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29811_ (.CLK(clknet_leaf_190_clk),
    .D(_00463_),
    .Q(\cpuregs[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29812_ (.CLK(clknet_leaf_188_clk),
    .D(_00464_),
    .Q(\cpuregs[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29813_ (.CLK(clknet_leaf_135_clk),
    .D(_00465_),
    .Q(\cpuregs[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29814_ (.CLK(clknet_leaf_145_clk),
    .D(_00466_),
    .Q(\cpuregs[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29815_ (.CLK(clknet_leaf_146_clk),
    .D(_00467_),
    .Q(\cpuregs[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29816_ (.CLK(clknet_leaf_136_clk),
    .D(_00468_),
    .Q(\cpuregs[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29817_ (.CLK(clknet_leaf_136_clk),
    .D(_00469_),
    .Q(\cpuregs[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29818_ (.CLK(clknet_leaf_134_clk),
    .D(_00470_),
    .Q(\cpuregs[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29819_ (.CLK(clknet_leaf_143_clk),
    .D(_00471_),
    .Q(\cpuregs[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29820_ (.CLK(clknet_leaf_147_clk),
    .D(_00472_),
    .Q(\cpuregs[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29821_ (.CLK(clknet_leaf_143_clk),
    .D(_00473_),
    .Q(\cpuregs[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29822_ (.CLK(clknet_leaf_147_clk),
    .D(_00474_),
    .Q(\cpuregs[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29823_ (.CLK(clknet_leaf_147_clk),
    .D(_00475_),
    .Q(\cpuregs[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29824_ (.CLK(clknet_leaf_143_clk),
    .D(_00476_),
    .Q(\cpuregs[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29825_ (.CLK(clknet_leaf_129_clk),
    .D(_00477_),
    .Q(\cpuregs[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29826_ (.CLK(clknet_leaf_125_clk),
    .D(_00478_),
    .Q(\cpuregs[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29827_ (.CLK(clknet_leaf_117_clk),
    .D(_00479_),
    .Q(\cpuregs[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29828_ (.CLK(clknet_leaf_128_clk),
    .D(_00480_),
    .Q(\cpuregs[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29829_ (.CLK(clknet_leaf_125_clk),
    .D(_00481_),
    .Q(\cpuregs[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29830_ (.CLK(clknet_leaf_117_clk),
    .D(_00482_),
    .Q(\cpuregs[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29831_ (.CLK(clknet_leaf_134_clk),
    .D(_00483_),
    .Q(\cpuregs[13][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29832_ (.CLK(clknet_leaf_146_clk),
    .D(_00484_),
    .Q(\cpuregs[13][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29833_ (.CLK(clknet_leaf_187_clk),
    .D(_00485_),
    .Q(\cpuregs[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29834_ (.CLK(clknet_leaf_178_clk),
    .D(_00486_),
    .Q(\cpuregs[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29835_ (.CLK(clknet_leaf_178_clk),
    .D(_00487_),
    .Q(\cpuregs[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29836_ (.CLK(clknet_leaf_188_clk),
    .D(_00488_),
    .Q(\cpuregs[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29837_ (.CLK(clknet_leaf_178_clk),
    .D(_00489_),
    .Q(\cpuregs[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29838_ (.CLK(clknet_leaf_187_clk),
    .D(_00490_),
    .Q(\cpuregs[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29839_ (.CLK(clknet_leaf_183_clk),
    .D(_00491_),
    .Q(\cpuregs[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29840_ (.CLK(clknet_leaf_193_clk),
    .D(_00492_),
    .Q(\cpuregs[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29841_ (.CLK(clknet_leaf_191_clk),
    .D(_00493_),
    .Q(\cpuregs[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29842_ (.CLK(clknet_leaf_152_clk),
    .D(_00494_),
    .Q(\cpuregs[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29843_ (.CLK(clknet_leaf_194_clk),
    .D(_00495_),
    .Q(\cpuregs[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29844_ (.CLK(clknet_leaf_188_clk),
    .D(_00496_),
    .Q(\cpuregs[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29845_ (.CLK(clknet_leaf_135_clk),
    .D(_00497_),
    .Q(\cpuregs[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29846_ (.CLK(clknet_leaf_135_clk),
    .D(_00498_),
    .Q(\cpuregs[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29847_ (.CLK(clknet_leaf_135_clk),
    .D(_00499_),
    .Q(\cpuregs[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29848_ (.CLK(clknet_leaf_135_clk),
    .D(_00500_),
    .Q(\cpuregs[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29849_ (.CLK(clknet_leaf_134_clk),
    .D(_00501_),
    .Q(\cpuregs[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29850_ (.CLK(clknet_leaf_134_clk),
    .D(_00502_),
    .Q(\cpuregs[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29851_ (.CLK(clknet_leaf_152_clk),
    .D(_00503_),
    .Q(\cpuregs[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29852_ (.CLK(clknet_leaf_152_clk),
    .D(_00504_),
    .Q(\cpuregs[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29853_ (.CLK(clknet_leaf_150_clk),
    .D(_00505_),
    .Q(\cpuregs[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29854_ (.CLK(clknet_leaf_152_clk),
    .D(_00506_),
    .Q(\cpuregs[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29855_ (.CLK(clknet_leaf_152_clk),
    .D(_00507_),
    .Q(\cpuregs[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29856_ (.CLK(clknet_leaf_152_clk),
    .D(_00508_),
    .Q(\cpuregs[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29857_ (.CLK(clknet_leaf_129_clk),
    .D(_00509_),
    .Q(\cpuregs[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29858_ (.CLK(clknet_leaf_138_clk),
    .D(_00510_),
    .Q(\cpuregs[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29859_ (.CLK(clknet_leaf_128_clk),
    .D(_00511_),
    .Q(\cpuregs[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29860_ (.CLK(clknet_leaf_128_clk),
    .D(_00512_),
    .Q(\cpuregs[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29861_ (.CLK(clknet_leaf_125_clk),
    .D(_00513_),
    .Q(\cpuregs[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29862_ (.CLK(clknet_leaf_128_clk),
    .D(_00514_),
    .Q(\cpuregs[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29863_ (.CLK(clknet_leaf_132_clk),
    .D(_00515_),
    .Q(\cpuregs[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29864_ (.CLK(clknet_leaf_146_clk),
    .D(_00516_),
    .Q(\cpuregs[14][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29865_ (.CLK(clknet_leaf_49_clk),
    .D(_00047_),
    .Q(\mem_wordsize[0] ));
 sky130_fd_sc_hd__dfxtp_1 _29866_ (.CLK(clknet_leaf_49_clk),
    .D(_00048_),
    .Q(\mem_wordsize[1] ));
 sky130_fd_sc_hd__dfxtp_2 _29867_ (.CLK(clknet_leaf_49_clk),
    .D(_00049_),
    .Q(\mem_wordsize[2] ));
 sky130_fd_sc_hd__dfxtp_1 _29868_ (.CLK(clknet_leaf_187_clk),
    .D(_00517_),
    .Q(\cpuregs[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29869_ (.CLK(clknet_leaf_178_clk),
    .D(_00518_),
    .Q(\cpuregs[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29870_ (.CLK(clknet_leaf_178_clk),
    .D(_00519_),
    .Q(\cpuregs[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29871_ (.CLK(clknet_leaf_188_clk),
    .D(_00520_),
    .Q(\cpuregs[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29872_ (.CLK(clknet_leaf_179_clk),
    .D(_00521_),
    .Q(\cpuregs[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29873_ (.CLK(clknet_leaf_158_clk),
    .D(_00522_),
    .Q(\cpuregs[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29874_ (.CLK(clknet_leaf_189_clk),
    .D(_00523_),
    .Q(\cpuregs[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29875_ (.CLK(clknet_leaf_193_clk),
    .D(_00524_),
    .Q(\cpuregs[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29876_ (.CLK(clknet_leaf_192_clk),
    .D(_00525_),
    .Q(\cpuregs[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29877_ (.CLK(clknet_leaf_192_clk),
    .D(_00526_),
    .Q(\cpuregs[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29878_ (.CLK(clknet_leaf_193_clk),
    .D(_00527_),
    .Q(\cpuregs[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29879_ (.CLK(clknet_leaf_189_clk),
    .D(_00528_),
    .Q(\cpuregs[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29880_ (.CLK(clknet_leaf_135_clk),
    .D(_00529_),
    .Q(\cpuregs[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29881_ (.CLK(clknet_leaf_135_clk),
    .D(_00530_),
    .Q(\cpuregs[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29882_ (.CLK(clknet_leaf_146_clk),
    .D(_00531_),
    .Q(\cpuregs[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29883_ (.CLK(clknet_leaf_135_clk),
    .D(_00532_),
    .Q(\cpuregs[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29884_ (.CLK(clknet_leaf_135_clk),
    .D(_00533_),
    .Q(\cpuregs[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29885_ (.CLK(clknet_leaf_135_clk),
    .D(_00534_),
    .Q(\cpuregs[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29886_ (.CLK(clknet_leaf_152_clk),
    .D(_00535_),
    .Q(\cpuregs[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29887_ (.CLK(clknet_leaf_152_clk),
    .D(_00536_),
    .Q(\cpuregs[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29888_ (.CLK(clknet_leaf_151_clk),
    .D(_00537_),
    .Q(\cpuregs[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29889_ (.CLK(clknet_leaf_152_clk),
    .D(_00538_),
    .Q(\cpuregs[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29890_ (.CLK(clknet_leaf_152_clk),
    .D(_00539_),
    .Q(\cpuregs[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29891_ (.CLK(clknet_leaf_152_clk),
    .D(_00540_),
    .Q(\cpuregs[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29892_ (.CLK(clknet_leaf_130_clk),
    .D(_00541_),
    .Q(\cpuregs[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29893_ (.CLK(clknet_leaf_133_clk),
    .D(_00542_),
    .Q(\cpuregs[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29894_ (.CLK(clknet_leaf_128_clk),
    .D(_00543_),
    .Q(\cpuregs[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29895_ (.CLK(clknet_leaf_128_clk),
    .D(_00544_),
    .Q(\cpuregs[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29896_ (.CLK(clknet_leaf_125_clk),
    .D(_00545_),
    .Q(\cpuregs[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29897_ (.CLK(clknet_leaf_127_clk),
    .D(_00546_),
    .Q(\cpuregs[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29898_ (.CLK(clknet_leaf_132_clk),
    .D(_00547_),
    .Q(\cpuregs[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29899_ (.CLK(clknet_leaf_147_clk),
    .D(_00548_),
    .Q(\cpuregs[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29900_ (.CLK(clknet_leaf_167_clk),
    .D(_00549_),
    .Q(\cpuregs[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29901_ (.CLK(clknet_leaf_174_clk),
    .D(_00550_),
    .Q(\cpuregs[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29902_ (.CLK(clknet_leaf_94_clk),
    .D(_00551_),
    .Q(\cpuregs[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29903_ (.CLK(clknet_leaf_97_clk),
    .D(_00552_),
    .Q(\cpuregs[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29904_ (.CLK(clknet_leaf_98_clk),
    .D(_00553_),
    .Q(\cpuregs[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29905_ (.CLK(clknet_leaf_97_clk),
    .D(_00554_),
    .Q(\cpuregs[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29906_ (.CLK(clknet_leaf_173_clk),
    .D(_00555_),
    .Q(\cpuregs[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29907_ (.CLK(clknet_leaf_99_clk),
    .D(_00556_),
    .Q(\cpuregs[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29908_ (.CLK(clknet_leaf_99_clk),
    .D(_00557_),
    .Q(\cpuregs[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29909_ (.CLK(clknet_leaf_168_clk),
    .D(_00558_),
    .Q(\cpuregs[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29910_ (.CLK(clknet_leaf_99_clk),
    .D(_00559_),
    .Q(\cpuregs[16][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29911_ (.CLK(clknet_leaf_167_clk),
    .D(_00560_),
    .Q(\cpuregs[16][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29912_ (.CLK(clknet_leaf_105_clk),
    .D(_00561_),
    .Q(\cpuregs[16][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29913_ (.CLK(clknet_leaf_105_clk),
    .D(_00562_),
    .Q(\cpuregs[16][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29914_ (.CLK(clknet_leaf_97_clk),
    .D(_00563_),
    .Q(\cpuregs[16][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29915_ (.CLK(clknet_leaf_102_clk),
    .D(_00564_),
    .Q(\cpuregs[16][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29916_ (.CLK(clknet_leaf_102_clk),
    .D(_00565_),
    .Q(\cpuregs[16][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29917_ (.CLK(clknet_leaf_105_clk),
    .D(_00566_),
    .Q(\cpuregs[16][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29918_ (.CLK(clknet_leaf_166_clk),
    .D(_00567_),
    .Q(\cpuregs[16][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29919_ (.CLK(clknet_leaf_165_clk),
    .D(_00568_),
    .Q(\cpuregs[16][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29920_ (.CLK(clknet_leaf_165_clk),
    .D(_00569_),
    .Q(\cpuregs[16][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29921_ (.CLK(clknet_leaf_165_clk),
    .D(_00570_),
    .Q(\cpuregs[16][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29922_ (.CLK(clknet_leaf_164_clk),
    .D(_00571_),
    .Q(\cpuregs[16][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29923_ (.CLK(clknet_leaf_98_clk),
    .D(_00572_),
    .Q(\cpuregs[16][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29924_ (.CLK(clknet_leaf_115_clk),
    .D(_00573_),
    .Q(\cpuregs[16][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29925_ (.CLK(clknet_leaf_120_clk),
    .D(_00574_),
    .Q(\cpuregs[16][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29926_ (.CLK(clknet_leaf_104_clk),
    .D(_00575_),
    .Q(\cpuregs[16][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29927_ (.CLK(clknet_leaf_114_clk),
    .D(_00576_),
    .Q(\cpuregs[16][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29928_ (.CLK(clknet_leaf_120_clk),
    .D(_00577_),
    .Q(\cpuregs[16][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29929_ (.CLK(clknet_leaf_114_clk),
    .D(_00578_),
    .Q(\cpuregs[16][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29930_ (.CLK(clknet_leaf_103_clk),
    .D(_00579_),
    .Q(\cpuregs[16][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29931_ (.CLK(clknet_leaf_97_clk),
    .D(_00580_),
    .Q(\cpuregs[16][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29932_ (.CLK(clknet_leaf_98_clk),
    .D(_00581_),
    .Q(\cpuregs[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29933_ (.CLK(clknet_leaf_173_clk),
    .D(_00582_),
    .Q(\cpuregs[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29934_ (.CLK(clknet_leaf_94_clk),
    .D(_00583_),
    .Q(\cpuregs[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29935_ (.CLK(clknet_leaf_97_clk),
    .D(_00584_),
    .Q(\cpuregs[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _29936_ (.CLK(clknet_leaf_98_clk),
    .D(_00585_),
    .Q(\cpuregs[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _29937_ (.CLK(clknet_leaf_97_clk),
    .D(_00586_),
    .Q(\cpuregs[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _29938_ (.CLK(clknet_leaf_167_clk),
    .D(_00587_),
    .Q(\cpuregs[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _29939_ (.CLK(clknet_leaf_99_clk),
    .D(_00588_),
    .Q(\cpuregs[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _29940_ (.CLK(clknet_leaf_99_clk),
    .D(_00589_),
    .Q(\cpuregs[17][8] ));
 sky130_fd_sc_hd__dfxtp_1 _29941_ (.CLK(clknet_leaf_168_clk),
    .D(_00590_),
    .Q(\cpuregs[17][9] ));
 sky130_fd_sc_hd__dfxtp_1 _29942_ (.CLK(clknet_leaf_99_clk),
    .D(_00591_),
    .Q(\cpuregs[17][10] ));
 sky130_fd_sc_hd__dfxtp_1 _29943_ (.CLK(clknet_leaf_167_clk),
    .D(_00592_),
    .Q(\cpuregs[17][11] ));
 sky130_fd_sc_hd__dfxtp_1 _29944_ (.CLK(clknet_leaf_105_clk),
    .D(_00593_),
    .Q(\cpuregs[17][12] ));
 sky130_fd_sc_hd__dfxtp_1 _29945_ (.CLK(clknet_leaf_105_clk),
    .D(_00594_),
    .Q(\cpuregs[17][13] ));
 sky130_fd_sc_hd__dfxtp_1 _29946_ (.CLK(clknet_leaf_97_clk),
    .D(_00595_),
    .Q(\cpuregs[17][14] ));
 sky130_fd_sc_hd__dfxtp_1 _29947_ (.CLK(clknet_leaf_99_clk),
    .D(_00596_),
    .Q(\cpuregs[17][15] ));
 sky130_fd_sc_hd__dfxtp_1 _29948_ (.CLK(clknet_leaf_102_clk),
    .D(_00597_),
    .Q(\cpuregs[17][16] ));
 sky130_fd_sc_hd__dfxtp_1 _29949_ (.CLK(clknet_leaf_104_clk),
    .D(_00598_),
    .Q(\cpuregs[17][17] ));
 sky130_fd_sc_hd__dfxtp_1 _29950_ (.CLK(clknet_leaf_166_clk),
    .D(_00599_),
    .Q(\cpuregs[17][18] ));
 sky130_fd_sc_hd__dfxtp_1 _29951_ (.CLK(clknet_leaf_163_clk),
    .D(_00600_),
    .Q(\cpuregs[17][19] ));
 sky130_fd_sc_hd__dfxtp_1 _29952_ (.CLK(clknet_leaf_165_clk),
    .D(_00601_),
    .Q(\cpuregs[17][20] ));
 sky130_fd_sc_hd__dfxtp_1 _29953_ (.CLK(clknet_leaf_165_clk),
    .D(_00602_),
    .Q(\cpuregs[17][21] ));
 sky130_fd_sc_hd__dfxtp_1 _29954_ (.CLK(clknet_leaf_165_clk),
    .D(_00603_),
    .Q(\cpuregs[17][22] ));
 sky130_fd_sc_hd__dfxtp_1 _29955_ (.CLK(clknet_leaf_166_clk),
    .D(_00604_),
    .Q(\cpuregs[17][23] ));
 sky130_fd_sc_hd__dfxtp_1 _29956_ (.CLK(clknet_leaf_120_clk),
    .D(_00605_),
    .Q(\cpuregs[17][24] ));
 sky130_fd_sc_hd__dfxtp_1 _29957_ (.CLK(clknet_leaf_120_clk),
    .D(_00606_),
    .Q(\cpuregs[17][25] ));
 sky130_fd_sc_hd__dfxtp_1 _29958_ (.CLK(clknet_leaf_104_clk),
    .D(_00607_),
    .Q(\cpuregs[17][26] ));
 sky130_fd_sc_hd__dfxtp_1 _29959_ (.CLK(clknet_leaf_115_clk),
    .D(_00608_),
    .Q(\cpuregs[17][27] ));
 sky130_fd_sc_hd__dfxtp_1 _29960_ (.CLK(clknet_leaf_121_clk),
    .D(_00609_),
    .Q(\cpuregs[17][28] ));
 sky130_fd_sc_hd__dfxtp_1 _29961_ (.CLK(clknet_leaf_115_clk),
    .D(_00610_),
    .Q(\cpuregs[17][29] ));
 sky130_fd_sc_hd__dfxtp_1 _29962_ (.CLK(clknet_leaf_121_clk),
    .D(_00611_),
    .Q(\cpuregs[17][30] ));
 sky130_fd_sc_hd__dfxtp_1 _29963_ (.CLK(clknet_leaf_97_clk),
    .D(_00612_),
    .Q(\cpuregs[17][31] ));
 sky130_fd_sc_hd__dfxtp_1 _29964_ (.CLK(clknet_leaf_66_clk),
    .D(_00613_),
    .Q(\mem_rdata_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _29965_ (.CLK(clknet_leaf_67_clk),
    .D(_00614_),
    .Q(\mem_rdata_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _29966_ (.CLK(clknet_leaf_67_clk),
    .D(_00615_),
    .Q(\mem_rdata_q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _29967_ (.CLK(clknet_leaf_86_clk),
    .D(_00616_),
    .Q(\mem_rdata_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _29968_ (.CLK(clknet_leaf_86_clk),
    .D(_00617_),
    .Q(\mem_rdata_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _29969_ (.CLK(clknet_leaf_64_clk),
    .D(_00618_),
    .Q(\mem_rdata_q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _29970_ (.CLK(clknet_leaf_64_clk),
    .D(_00619_),
    .Q(\mem_rdata_q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _29971_ (.CLK(clknet_leaf_84_clk),
    .D(_00620_),
    .Q(\mem_rdata_q[7] ));
 sky130_fd_sc_hd__dfxtp_2 _29972_ (.CLK(clknet_leaf_84_clk),
    .D(_00621_),
    .Q(\mem_rdata_q[8] ));
 sky130_fd_sc_hd__dfxtp_2 _29973_ (.CLK(clknet_leaf_83_clk),
    .D(_00622_),
    .Q(\mem_rdata_q[9] ));
 sky130_fd_sc_hd__dfxtp_2 _29974_ (.CLK(clknet_leaf_67_clk),
    .D(_00623_),
    .Q(\mem_rdata_q[10] ));
 sky130_fd_sc_hd__dfxtp_2 _29975_ (.CLK(clknet_leaf_87_clk),
    .D(_00624_),
    .Q(\mem_rdata_q[11] ));
 sky130_fd_sc_hd__dfxtp_2 _29976_ (.CLK(clknet_leaf_33_clk),
    .D(_00625_),
    .Q(\mem_rdata_q[12] ));
 sky130_fd_sc_hd__dfxtp_1 _29977_ (.CLK(clknet_leaf_32_clk),
    .D(_00626_),
    .Q(\mem_rdata_q[13] ));
 sky130_fd_sc_hd__dfxtp_2 _29978_ (.CLK(clknet_leaf_32_clk),
    .D(_00627_),
    .Q(\mem_rdata_q[14] ));
 sky130_fd_sc_hd__dfxtp_2 _29979_ (.CLK(clknet_leaf_30_clk),
    .D(_00628_),
    .Q(\mem_rdata_q[15] ));
 sky130_fd_sc_hd__dfxtp_2 _29980_ (.CLK(clknet_leaf_88_clk),
    .D(_00629_),
    .Q(\mem_rdata_q[16] ));
 sky130_fd_sc_hd__dfxtp_2 _29981_ (.CLK(clknet_leaf_88_clk),
    .D(_00630_),
    .Q(\mem_rdata_q[17] ));
 sky130_fd_sc_hd__dfxtp_2 _29982_ (.CLK(clknet_leaf_88_clk),
    .D(_00631_),
    .Q(\mem_rdata_q[18] ));
 sky130_fd_sc_hd__dfxtp_2 _29983_ (.CLK(clknet_leaf_88_clk),
    .D(_00632_),
    .Q(\mem_rdata_q[19] ));
 sky130_fd_sc_hd__dfxtp_4 _29984_ (.CLK(clknet_leaf_30_clk),
    .D(_00633_),
    .Q(\mem_rdata_q[20] ));
 sky130_fd_sc_hd__dfxtp_2 _29985_ (.CLK(clknet_leaf_31_clk),
    .D(_00634_),
    .Q(\mem_rdata_q[21] ));
 sky130_fd_sc_hd__dfxtp_2 _29986_ (.CLK(clknet_leaf_31_clk),
    .D(_00635_),
    .Q(\mem_rdata_q[22] ));
 sky130_fd_sc_hd__dfxtp_2 _29987_ (.CLK(clknet_leaf_31_clk),
    .D(_00636_),
    .Q(\mem_rdata_q[23] ));
 sky130_fd_sc_hd__dfxtp_2 _29988_ (.CLK(clknet_leaf_30_clk),
    .D(_00637_),
    .Q(\mem_rdata_q[24] ));
 sky130_fd_sc_hd__dfxtp_1 _29989_ (.CLK(clknet_leaf_87_clk),
    .D(_00638_),
    .Q(\mem_rdata_q[25] ));
 sky130_fd_sc_hd__dfxtp_1 _29990_ (.CLK(clknet_leaf_30_clk),
    .D(_00639_),
    .Q(\mem_rdata_q[26] ));
 sky130_fd_sc_hd__dfxtp_1 _29991_ (.CLK(clknet_leaf_87_clk),
    .D(_00640_),
    .Q(\mem_rdata_q[27] ));
 sky130_fd_sc_hd__dfxtp_2 _29992_ (.CLK(clknet_leaf_29_clk),
    .D(_00641_),
    .Q(\mem_rdata_q[28] ));
 sky130_fd_sc_hd__dfxtp_1 _29993_ (.CLK(clknet_leaf_31_clk),
    .D(_00642_),
    .Q(\mem_rdata_q[29] ));
 sky130_fd_sc_hd__dfxtp_1 _29994_ (.CLK(clknet_leaf_31_clk),
    .D(_00643_),
    .Q(\mem_rdata_q[30] ));
 sky130_fd_sc_hd__dfxtp_1 _29995_ (.CLK(clknet_leaf_29_clk),
    .D(_00644_),
    .Q(\mem_rdata_q[31] ));
 sky130_fd_sc_hd__dfxtp_1 _29996_ (.CLK(clknet_leaf_167_clk),
    .D(_00645_),
    .Q(\cpuregs[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _29997_ (.CLK(clknet_leaf_173_clk),
    .D(_00646_),
    .Q(\cpuregs[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _29998_ (.CLK(clknet_leaf_173_clk),
    .D(_00647_),
    .Q(\cpuregs[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _29999_ (.CLK(clknet_leaf_98_clk),
    .D(_00648_),
    .Q(\cpuregs[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30000_ (.CLK(clknet_leaf_166_clk),
    .D(_00649_),
    .Q(\cpuregs[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30001_ (.CLK(clknet_leaf_98_clk),
    .D(_00650_),
    .Q(\cpuregs[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30002_ (.CLK(clknet_leaf_167_clk),
    .D(_00651_),
    .Q(\cpuregs[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30003_ (.CLK(clknet_leaf_166_clk),
    .D(_00652_),
    .Q(\cpuregs[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30004_ (.CLK(clknet_leaf_166_clk),
    .D(_00653_),
    .Q(\cpuregs[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30005_ (.CLK(clknet_leaf_168_clk),
    .D(_00654_),
    .Q(\cpuregs[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30006_ (.CLK(clknet_leaf_98_clk),
    .D(_00655_),
    .Q(\cpuregs[18][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30007_ (.CLK(clknet_leaf_168_clk),
    .D(_00656_),
    .Q(\cpuregs[18][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30008_ (.CLK(clknet_leaf_102_clk),
    .D(_00657_),
    .Q(\cpuregs[18][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30009_ (.CLK(clknet_leaf_102_clk),
    .D(_00658_),
    .Q(\cpuregs[18][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30010_ (.CLK(clknet_leaf_102_clk),
    .D(_00659_),
    .Q(\cpuregs[18][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30011_ (.CLK(clknet_leaf_101_clk),
    .D(_00660_),
    .Q(\cpuregs[18][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30012_ (.CLK(clknet_leaf_102_clk),
    .D(_00661_),
    .Q(\cpuregs[18][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30013_ (.CLK(clknet_leaf_103_clk),
    .D(_00662_),
    .Q(\cpuregs[18][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30014_ (.CLK(clknet_leaf_165_clk),
    .D(_00663_),
    .Q(\cpuregs[18][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30015_ (.CLK(clknet_leaf_163_clk),
    .D(_00664_),
    .Q(\cpuregs[18][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30016_ (.CLK(clknet_leaf_164_clk),
    .D(_00665_),
    .Q(\cpuregs[18][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30017_ (.CLK(clknet_leaf_163_clk),
    .D(_00666_),
    .Q(\cpuregs[18][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30018_ (.CLK(clknet_leaf_163_clk),
    .D(_00667_),
    .Q(\cpuregs[18][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30019_ (.CLK(clknet_leaf_162_clk),
    .D(_00668_),
    .Q(\cpuregs[18][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30020_ (.CLK(clknet_leaf_116_clk),
    .D(_00669_),
    .Q(\cpuregs[18][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30021_ (.CLK(clknet_leaf_120_clk),
    .D(_00670_),
    .Q(\cpuregs[18][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30022_ (.CLK(clknet_leaf_115_clk),
    .D(_00671_),
    .Q(\cpuregs[18][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30023_ (.CLK(clknet_leaf_115_clk),
    .D(_00672_),
    .Q(\cpuregs[18][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30024_ (.CLK(clknet_leaf_121_clk),
    .D(_00673_),
    .Q(\cpuregs[18][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30025_ (.CLK(clknet_leaf_116_clk),
    .D(_00674_),
    .Q(\cpuregs[18][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30026_ (.CLK(clknet_leaf_121_clk),
    .D(_00675_),
    .Q(\cpuregs[18][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30027_ (.CLK(clknet_leaf_99_clk),
    .D(_00676_),
    .Q(\cpuregs[18][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30028_ (.CLK(clknet_leaf_159_clk),
    .D(_00677_),
    .Q(\cpuregs[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30029_ (.CLK(clknet_leaf_172_clk),
    .D(_00678_),
    .Q(\cpuregs[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30030_ (.CLK(clknet_leaf_171_clk),
    .D(_00679_),
    .Q(\cpuregs[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30031_ (.CLK(clknet_leaf_168_clk),
    .D(_00680_),
    .Q(\cpuregs[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30032_ (.CLK(clknet_leaf_169_clk),
    .D(_00681_),
    .Q(\cpuregs[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30033_ (.CLK(clknet_leaf_169_clk),
    .D(_00682_),
    .Q(\cpuregs[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30034_ (.CLK(clknet_leaf_186_clk),
    .D(_00683_),
    .Q(\cpuregs[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30035_ (.CLK(clknet_leaf_192_clk),
    .D(_00684_),
    .Q(\cpuregs[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30036_ (.CLK(clknet_leaf_152_clk),
    .D(_00685_),
    .Q(\cpuregs[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30037_ (.CLK(clknet_leaf_153_clk),
    .D(_00686_),
    .Q(\cpuregs[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30038_ (.CLK(clknet_leaf_189_clk),
    .D(_00687_),
    .Q(\cpuregs[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30039_ (.CLK(clknet_leaf_156_clk),
    .D(_00688_),
    .Q(\cpuregs[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30040_ (.CLK(clknet_leaf_136_clk),
    .D(_00689_),
    .Q(\cpuregs[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30041_ (.CLK(clknet_leaf_123_clk),
    .D(_00690_),
    .Q(\cpuregs[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30042_ (.CLK(clknet_leaf_164_clk),
    .D(_00691_),
    .Q(\cpuregs[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30043_ (.CLK(clknet_leaf_140_clk),
    .D(_00692_),
    .Q(\cpuregs[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30044_ (.CLK(clknet_leaf_137_clk),
    .D(_00693_),
    .Q(\cpuregs[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30045_ (.CLK(clknet_leaf_124_clk),
    .D(_00694_),
    .Q(\cpuregs[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30046_ (.CLK(clknet_leaf_143_clk),
    .D(_00695_),
    .Q(\cpuregs[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30047_ (.CLK(clknet_leaf_143_clk),
    .D(_00696_),
    .Q(\cpuregs[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30048_ (.CLK(clknet_leaf_143_clk),
    .D(_00697_),
    .Q(\cpuregs[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30049_ (.CLK(clknet_leaf_142_clk),
    .D(_00698_),
    .Q(\cpuregs[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30050_ (.CLK(clknet_leaf_144_clk),
    .D(_00699_),
    .Q(\cpuregs[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30051_ (.CLK(clknet_leaf_161_clk),
    .D(_00700_),
    .Q(\cpuregs[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30052_ (.CLK(clknet_leaf_129_clk),
    .D(_00701_),
    .Q(\cpuregs[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30053_ (.CLK(clknet_leaf_125_clk),
    .D(_00702_),
    .Q(\cpuregs[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30054_ (.CLK(clknet_leaf_116_clk),
    .D(_00703_),
    .Q(\cpuregs[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30055_ (.CLK(clknet_leaf_119_clk),
    .D(_00704_),
    .Q(\cpuregs[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30056_ (.CLK(clknet_leaf_126_clk),
    .D(_00705_),
    .Q(\cpuregs[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30057_ (.CLK(clknet_leaf_116_clk),
    .D(_00706_),
    .Q(\cpuregs[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30058_ (.CLK(clknet_leaf_134_clk),
    .D(_00707_),
    .Q(\cpuregs[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30059_ (.CLK(clknet_leaf_146_clk),
    .D(_00708_),
    .Q(\cpuregs[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30060_ (.CLK(clknet_leaf_213_clk),
    .D(_00709_),
    .Q(\genblk1.pcpi_mul.rs1[0] ));
 sky130_fd_sc_hd__dfxtp_2 _30061_ (.CLK(clknet_leaf_213_clk),
    .D(_00710_),
    .Q(\genblk1.pcpi_mul.rs1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _30062_ (.CLK(clknet_leaf_213_clk),
    .D(_00711_),
    .Q(\genblk1.pcpi_mul.rs1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30063_ (.CLK(clknet_leaf_213_clk),
    .D(_00712_),
    .Q(\genblk1.pcpi_mul.rs1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30064_ (.CLK(clknet_leaf_217_clk),
    .D(_00713_),
    .Q(\genblk1.pcpi_mul.rs1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _30065_ (.CLK(clknet_leaf_217_clk),
    .D(_00714_),
    .Q(\genblk1.pcpi_mul.rs1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _30066_ (.CLK(clknet_5_4__leaf_clk),
    .D(_00715_),
    .Q(\genblk1.pcpi_mul.rs1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _30067_ (.CLK(clknet_leaf_218_clk),
    .D(_00716_),
    .Q(\genblk1.pcpi_mul.rs1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _30068_ (.CLK(clknet_leaf_219_clk),
    .D(_00717_),
    .Q(\genblk1.pcpi_mul.rs1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _30069_ (.CLK(clknet_leaf_219_clk),
    .D(_00718_),
    .Q(\genblk1.pcpi_mul.rs1[9] ));
 sky130_fd_sc_hd__dfxtp_2 _30070_ (.CLK(clknet_leaf_224_clk),
    .D(_00719_),
    .Q(\genblk1.pcpi_mul.rs1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _30071_ (.CLK(clknet_leaf_224_clk),
    .D(_00720_),
    .Q(\genblk1.pcpi_mul.rs1[11] ));
 sky130_fd_sc_hd__dfxtp_2 _30072_ (.CLK(clknet_leaf_224_clk),
    .D(_00721_),
    .Q(\genblk1.pcpi_mul.rs1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _30073_ (.CLK(clknet_leaf_0_clk),
    .D(_00722_),
    .Q(\genblk1.pcpi_mul.rs1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _30074_ (.CLK(clknet_leaf_224_clk),
    .D(_00723_),
    .Q(\genblk1.pcpi_mul.rs1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _30075_ (.CLK(clknet_leaf_224_clk),
    .D(_00724_),
    .Q(\genblk1.pcpi_mul.rs1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _30076_ (.CLK(clknet_5_1__leaf_clk),
    .D(_00725_),
    .Q(\genblk1.pcpi_mul.rs1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _30077_ (.CLK(clknet_leaf_221_clk),
    .D(_00726_),
    .Q(\genblk1.pcpi_mul.rs1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _30078_ (.CLK(clknet_leaf_221_clk),
    .D(_00727_),
    .Q(\genblk1.pcpi_mul.rs1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _30079_ (.CLK(clknet_leaf_221_clk),
    .D(_00728_),
    .Q(\genblk1.pcpi_mul.rs1[19] ));
 sky130_fd_sc_hd__dfxtp_2 _30080_ (.CLK(clknet_leaf_196_clk),
    .D(_00729_),
    .Q(\genblk1.pcpi_mul.rs1[20] ));
 sky130_fd_sc_hd__dfxtp_2 _30081_ (.CLK(clknet_leaf_196_clk),
    .D(_00730_),
    .Q(\genblk1.pcpi_mul.rs1[21] ));
 sky130_fd_sc_hd__dfxtp_2 _30082_ (.CLK(clknet_leaf_196_clk),
    .D(_00731_),
    .Q(\genblk1.pcpi_mul.rs1[22] ));
 sky130_fd_sc_hd__dfxtp_4 _30083_ (.CLK(clknet_leaf_196_clk),
    .D(_00732_),
    .Q(\genblk1.pcpi_mul.rs1[23] ));
 sky130_fd_sc_hd__dfxtp_2 _30084_ (.CLK(clknet_leaf_196_clk),
    .D(_00733_),
    .Q(\genblk1.pcpi_mul.rs1[24] ));
 sky130_fd_sc_hd__dfxtp_2 _30085_ (.CLK(clknet_leaf_197_clk),
    .D(_00734_),
    .Q(\genblk1.pcpi_mul.rs1[25] ));
 sky130_fd_sc_hd__dfxtp_4 _30086_ (.CLK(clknet_leaf_197_clk),
    .D(_00735_),
    .Q(\genblk1.pcpi_mul.rs1[26] ));
 sky130_fd_sc_hd__dfxtp_4 _30087_ (.CLK(clknet_leaf_204_clk),
    .D(_00736_),
    .Q(\genblk1.pcpi_mul.rs1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _30088_ (.CLK(clknet_leaf_198_clk),
    .D(_00737_),
    .Q(\genblk1.pcpi_mul.rs1[28] ));
 sky130_fd_sc_hd__dfxtp_2 _30089_ (.CLK(clknet_5_16__leaf_clk),
    .D(_00738_),
    .Q(\genblk1.pcpi_mul.rs1[29] ));
 sky130_fd_sc_hd__dfxtp_4 _30090_ (.CLK(clknet_leaf_204_clk),
    .D(_00739_),
    .Q(\genblk1.pcpi_mul.rs1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _30091_ (.CLK(clknet_leaf_198_clk),
    .D(_00740_),
    .Q(\genblk1.pcpi_mul.rs1[31] ));
 sky130_fd_sc_hd__dfxtp_2 _30092_ (.CLK(clknet_leaf_204_clk),
    .D(_00741_),
    .Q(\genblk1.pcpi_mul.rs2[0] ));
 sky130_fd_sc_hd__dfxtp_2 _30093_ (.CLK(clknet_leaf_204_clk),
    .D(_00742_),
    .Q(\genblk1.pcpi_mul.rs2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30094_ (.CLK(clknet_leaf_214_clk),
    .D(_00743_),
    .Q(\genblk1.pcpi_mul.rs2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30095_ (.CLK(clknet_leaf_214_clk),
    .D(_00744_),
    .Q(\genblk1.pcpi_mul.rs2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30096_ (.CLK(clknet_leaf_218_clk),
    .D(_00745_),
    .Q(\genblk1.pcpi_mul.rs2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _30097_ (.CLK(clknet_leaf_218_clk),
    .D(_00746_),
    .Q(\genblk1.pcpi_mul.rs2[5] ));
 sky130_fd_sc_hd__dfxtp_2 _30098_ (.CLK(clknet_leaf_214_clk),
    .D(_00747_),
    .Q(\genblk1.pcpi_mul.rs2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _30099_ (.CLK(clknet_leaf_218_clk),
    .D(_00748_),
    .Q(\genblk1.pcpi_mul.rs2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _30100_ (.CLK(clknet_leaf_218_clk),
    .D(_00749_),
    .Q(\genblk1.pcpi_mul.rs2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _30101_ (.CLK(clknet_leaf_218_clk),
    .D(_00750_),
    .Q(\genblk1.pcpi_mul.rs2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _30102_ (.CLK(clknet_leaf_224_clk),
    .D(_00751_),
    .Q(\genblk1.pcpi_mul.rs2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _30103_ (.CLK(clknet_leaf_218_clk),
    .D(_00752_),
    .Q(\genblk1.pcpi_mul.rs2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _30104_ (.CLK(clknet_leaf_224_clk),
    .D(_00753_),
    .Q(\genblk1.pcpi_mul.rs2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _30105_ (.CLK(clknet_leaf_224_clk),
    .D(_00754_),
    .Q(\genblk1.pcpi_mul.rs2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _30106_ (.CLK(clknet_leaf_0_clk),
    .D(_00755_),
    .Q(\genblk1.pcpi_mul.rs2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _30107_ (.CLK(clknet_leaf_225_clk),
    .D(_00756_),
    .Q(\genblk1.pcpi_mul.rs2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _30108_ (.CLK(clknet_leaf_16_clk),
    .D(_00757_),
    .Q(\genblk1.pcpi_mul.rs2[16] ));
 sky130_fd_sc_hd__dfxtp_2 _30109_ (.CLK(clknet_leaf_16_clk),
    .D(_00758_),
    .Q(\genblk1.pcpi_mul.rs2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _30110_ (.CLK(clknet_leaf_16_clk),
    .D(_00759_),
    .Q(\genblk1.pcpi_mul.rs2[18] ));
 sky130_fd_sc_hd__dfxtp_1 _30111_ (.CLK(clknet_leaf_16_clk),
    .D(_00760_),
    .Q(\genblk1.pcpi_mul.rs2[19] ));
 sky130_fd_sc_hd__dfxtp_1 _30112_ (.CLK(clknet_leaf_217_clk),
    .D(_00761_),
    .Q(\genblk1.pcpi_mul.rs2[20] ));
 sky130_fd_sc_hd__dfxtp_2 _30113_ (.CLK(clknet_leaf_214_clk),
    .D(_00762_),
    .Q(\genblk1.pcpi_mul.rs2[21] ));
 sky130_fd_sc_hd__dfxtp_1 _30114_ (.CLK(clknet_leaf_216_clk),
    .D(_00763_),
    .Q(\genblk1.pcpi_mul.rs2[22] ));
 sky130_fd_sc_hd__dfxtp_1 _30115_ (.CLK(clknet_leaf_216_clk),
    .D(_00764_),
    .Q(\genblk1.pcpi_mul.rs2[23] ));
 sky130_fd_sc_hd__dfxtp_1 _30116_ (.CLK(clknet_leaf_216_clk),
    .D(_00765_),
    .Q(\genblk1.pcpi_mul.rs2[24] ));
 sky130_fd_sc_hd__dfxtp_1 _30117_ (.CLK(clknet_leaf_216_clk),
    .D(_00766_),
    .Q(\genblk1.pcpi_mul.rs2[25] ));
 sky130_fd_sc_hd__dfxtp_1 _30118_ (.CLK(clknet_leaf_216_clk),
    .D(_00767_),
    .Q(\genblk1.pcpi_mul.rs2[26] ));
 sky130_fd_sc_hd__dfxtp_1 _30119_ (.CLK(clknet_leaf_216_clk),
    .D(_00768_),
    .Q(\genblk1.pcpi_mul.rs2[27] ));
 sky130_fd_sc_hd__dfxtp_1 _30120_ (.CLK(clknet_leaf_215_clk),
    .D(_00769_),
    .Q(\genblk1.pcpi_mul.rs2[28] ));
 sky130_fd_sc_hd__dfxtp_1 _30121_ (.CLK(clknet_leaf_216_clk),
    .D(_00770_),
    .Q(\genblk1.pcpi_mul.rs2[29] ));
 sky130_fd_sc_hd__dfxtp_1 _30122_ (.CLK(clknet_leaf_215_clk),
    .D(_00771_),
    .Q(\genblk1.pcpi_mul.rs2[30] ));
 sky130_fd_sc_hd__dfxtp_1 _30123_ (.CLK(clknet_leaf_215_clk),
    .D(_00772_),
    .Q(\genblk1.pcpi_mul.rs2[31] ));
 sky130_fd_sc_hd__dfxtp_1 _30124_ (.CLK(clknet_leaf_83_clk),
    .D(_00036_),
    .Q(\irq_pending[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30125_ (.CLK(clknet_leaf_50_clk),
    .D(_00773_),
    .Q(\genblk1.pcpi_mul.active[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30126_ (.CLK(clknet_leaf_64_clk),
    .D(_00774_),
    .Q(\genblk1.pcpi_mul.active[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30127_ (.CLK(clknet_leaf_83_clk),
    .D(_00775_),
    .Q(net331));
 sky130_fd_sc_hd__dfxtp_2 _30128_ (.CLK(clknet_leaf_108_clk),
    .D(_00776_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_1 _30129_ (.CLK(clknet_leaf_108_clk),
    .D(_00777_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_1 _30130_ (.CLK(clknet_leaf_108_clk),
    .D(_00778_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_1 _30131_ (.CLK(clknet_leaf_108_clk),
    .D(_00779_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_1 _30132_ (.CLK(clknet_leaf_108_clk),
    .D(_00780_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_1 _30133_ (.CLK(clknet_leaf_108_clk),
    .D(_00781_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_1 _30134_ (.CLK(clknet_leaf_109_clk),
    .D(_00782_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_1 _30135_ (.CLK(clknet_leaf_108_clk),
    .D(_00783_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_1 _30136_ (.CLK(clknet_leaf_109_clk),
    .D(_00784_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_1 _30137_ (.CLK(clknet_leaf_109_clk),
    .D(_00785_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_1 _30138_ (.CLK(clknet_leaf_105_clk),
    .D(_00786_),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_1 _30139_ (.CLK(clknet_leaf_105_clk),
    .D(_00787_),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_1 _30140_ (.CLK(clknet_leaf_106_clk),
    .D(_00788_),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_1 _30141_ (.CLK(clknet_leaf_106_clk),
    .D(_00789_),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_1 _30142_ (.CLK(clknet_leaf_105_clk),
    .D(_00790_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_1 _30143_ (.CLK(clknet_leaf_106_clk),
    .D(_00791_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_1 _30144_ (.CLK(clknet_leaf_106_clk),
    .D(_00792_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_1 _30145_ (.CLK(clknet_leaf_106_clk),
    .D(_00793_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_1 _30146_ (.CLK(clknet_leaf_96_clk),
    .D(_00794_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_1 _30147_ (.CLK(clknet_leaf_96_clk),
    .D(_00795_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_1 _30148_ (.CLK(clknet_leaf_96_clk),
    .D(_00796_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_1 _30149_ (.CLK(clknet_leaf_96_clk),
    .D(_00797_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_1 _30150_ (.CLK(clknet_leaf_96_clk),
    .D(_00798_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_1 _30151_ (.CLK(clknet_leaf_106_clk),
    .D(_00799_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_1 _30152_ (.CLK(clknet_leaf_106_clk),
    .D(_00800_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_2 _30153_ (.CLK(clknet_leaf_96_clk),
    .D(_00801_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_2 _30154_ (.CLK(clknet_leaf_106_clk),
    .D(_00802_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_1 _30155_ (.CLK(clknet_leaf_106_clk),
    .D(_00803_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_1 _30156_ (.CLK(clknet_leaf_107_clk),
    .D(_00804_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_1 _30157_ (.CLK(clknet_leaf_107_clk),
    .D(_00805_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_1 _30158_ (.CLK(clknet_leaf_107_clk),
    .D(_00806_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_1 _30159_ (.CLK(clknet_leaf_108_clk),
    .D(_00807_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_1 _30160_ (.CLK(clknet_leaf_83_clk),
    .D(_00808_),
    .Q(net332));
 sky130_fd_sc_hd__dfxtp_1 _30161_ (.CLK(clknet_leaf_73_clk),
    .D(_00809_),
    .Q(\count_instr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30162_ (.CLK(clknet_leaf_73_clk),
    .D(_00810_),
    .Q(\count_instr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30163_ (.CLK(clknet_leaf_73_clk),
    .D(_00811_),
    .Q(\count_instr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30164_ (.CLK(clknet_leaf_72_clk),
    .D(_00812_),
    .Q(\count_instr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30165_ (.CLK(clknet_leaf_71_clk),
    .D(_00813_),
    .Q(\count_instr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _30166_ (.CLK(clknet_leaf_71_clk),
    .D(_00814_),
    .Q(\count_instr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _30167_ (.CLK(clknet_leaf_72_clk),
    .D(_00815_),
    .Q(\count_instr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _30168_ (.CLK(clknet_leaf_68_clk),
    .D(_00816_),
    .Q(\count_instr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _30169_ (.CLK(clknet_leaf_68_clk),
    .D(_00817_),
    .Q(\count_instr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _30170_ (.CLK(clknet_leaf_68_clk),
    .D(_00818_),
    .Q(\count_instr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _30171_ (.CLK(clknet_leaf_60_clk),
    .D(_00819_),
    .Q(\count_instr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _30172_ (.CLK(clknet_leaf_60_clk),
    .D(_00820_),
    .Q(\count_instr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _30173_ (.CLK(clknet_leaf_61_clk),
    .D(_00821_),
    .Q(\count_instr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _30174_ (.CLK(clknet_leaf_61_clk),
    .D(_00822_),
    .Q(\count_instr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _30175_ (.CLK(clknet_leaf_61_clk),
    .D(_00823_),
    .Q(\count_instr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _30176_ (.CLK(clknet_leaf_63_clk),
    .D(_00824_),
    .Q(\count_instr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _30177_ (.CLK(clknet_leaf_63_clk),
    .D(_00825_),
    .Q(\count_instr[16] ));
 sky130_fd_sc_hd__dfxtp_1 _30178_ (.CLK(clknet_leaf_63_clk),
    .D(_00826_),
    .Q(\count_instr[17] ));
 sky130_fd_sc_hd__dfxtp_1 _30179_ (.CLK(clknet_leaf_61_clk),
    .D(_00827_),
    .Q(\count_instr[18] ));
 sky130_fd_sc_hd__dfxtp_1 _30180_ (.CLK(clknet_leaf_62_clk),
    .D(_00828_),
    .Q(\count_instr[19] ));
 sky130_fd_sc_hd__dfxtp_1 _30181_ (.CLK(clknet_leaf_62_clk),
    .D(_00829_),
    .Q(\count_instr[20] ));
 sky130_fd_sc_hd__dfxtp_1 _30182_ (.CLK(clknet_leaf_62_clk),
    .D(_00830_),
    .Q(\count_instr[21] ));
 sky130_fd_sc_hd__dfxtp_1 _30183_ (.CLK(clknet_leaf_56_clk),
    .D(_00831_),
    .Q(\count_instr[22] ));
 sky130_fd_sc_hd__dfxtp_1 _30184_ (.CLK(clknet_leaf_62_clk),
    .D(_00832_),
    .Q(\count_instr[23] ));
 sky130_fd_sc_hd__dfxtp_1 _30185_ (.CLK(clknet_leaf_61_clk),
    .D(_00833_),
    .Q(\count_instr[24] ));
 sky130_fd_sc_hd__dfxtp_1 _30186_ (.CLK(clknet_leaf_57_clk),
    .D(_00834_),
    .Q(\count_instr[25] ));
 sky130_fd_sc_hd__dfxtp_1 _30187_ (.CLK(clknet_leaf_58_clk),
    .D(_00835_),
    .Q(\count_instr[26] ));
 sky130_fd_sc_hd__dfxtp_1 _30188_ (.CLK(clknet_leaf_60_clk),
    .D(_00836_),
    .Q(\count_instr[27] ));
 sky130_fd_sc_hd__dfxtp_1 _30189_ (.CLK(clknet_leaf_58_clk),
    .D(_00837_),
    .Q(\count_instr[28] ));
 sky130_fd_sc_hd__dfxtp_1 _30190_ (.CLK(clknet_leaf_59_clk),
    .D(_00838_),
    .Q(\count_instr[29] ));
 sky130_fd_sc_hd__dfxtp_1 _30191_ (.CLK(clknet_leaf_59_clk),
    .D(_00839_),
    .Q(\count_instr[30] ));
 sky130_fd_sc_hd__dfxtp_1 _30192_ (.CLK(clknet_leaf_70_clk),
    .D(_00840_),
    .Q(\count_instr[31] ));
 sky130_fd_sc_hd__dfxtp_1 _30193_ (.CLK(clknet_leaf_70_clk),
    .D(_00841_),
    .Q(\count_instr[32] ));
 sky130_fd_sc_hd__dfxtp_1 _30194_ (.CLK(clknet_leaf_71_clk),
    .D(_00842_),
    .Q(\count_instr[33] ));
 sky130_fd_sc_hd__dfxtp_1 _30195_ (.CLK(clknet_leaf_70_clk),
    .D(_00843_),
    .Q(\count_instr[34] ));
 sky130_fd_sc_hd__dfxtp_1 _30196_ (.CLK(clknet_leaf_70_clk),
    .D(_00844_),
    .Q(\count_instr[35] ));
 sky130_fd_sc_hd__dfxtp_1 _30197_ (.CLK(clknet_leaf_68_clk),
    .D(_00845_),
    .Q(\count_instr[36] ));
 sky130_fd_sc_hd__dfxtp_1 _30198_ (.CLK(clknet_leaf_68_clk),
    .D(_00846_),
    .Q(\count_instr[37] ));
 sky130_fd_sc_hd__dfxtp_1 _30199_ (.CLK(clknet_leaf_70_clk),
    .D(_00847_),
    .Q(\count_instr[38] ));
 sky130_fd_sc_hd__dfxtp_1 _30200_ (.CLK(clknet_leaf_69_clk),
    .D(_00848_),
    .Q(\count_instr[39] ));
 sky130_fd_sc_hd__dfxtp_1 _30201_ (.CLK(clknet_leaf_69_clk),
    .D(_00849_),
    .Q(\count_instr[40] ));
 sky130_fd_sc_hd__dfxtp_1 _30202_ (.CLK(clknet_leaf_69_clk),
    .D(_00850_),
    .Q(\count_instr[41] ));
 sky130_fd_sc_hd__dfxtp_1 _30203_ (.CLK(clknet_leaf_60_clk),
    .D(_00851_),
    .Q(\count_instr[42] ));
 sky130_fd_sc_hd__dfxtp_1 _30204_ (.CLK(clknet_leaf_59_clk),
    .D(_00852_),
    .Q(\count_instr[43] ));
 sky130_fd_sc_hd__dfxtp_1 _30205_ (.CLK(clknet_leaf_59_clk),
    .D(_00853_),
    .Q(\count_instr[44] ));
 sky130_fd_sc_hd__dfxtp_1 _30206_ (.CLK(clknet_leaf_58_clk),
    .D(_00854_),
    .Q(\count_instr[45] ));
 sky130_fd_sc_hd__dfxtp_1 _30207_ (.CLK(clknet_leaf_58_clk),
    .D(_00855_),
    .Q(\count_instr[46] ));
 sky130_fd_sc_hd__dfxtp_1 _30208_ (.CLK(clknet_leaf_58_clk),
    .D(_00856_),
    .Q(\count_instr[47] ));
 sky130_fd_sc_hd__dfxtp_1 _30209_ (.CLK(clknet_leaf_58_clk),
    .D(_00857_),
    .Q(\count_instr[48] ));
 sky130_fd_sc_hd__dfxtp_1 _30210_ (.CLK(clknet_leaf_57_clk),
    .D(_00858_),
    .Q(\count_instr[49] ));
 sky130_fd_sc_hd__dfxtp_1 _30211_ (.CLK(clknet_leaf_55_clk),
    .D(_00859_),
    .Q(\count_instr[50] ));
 sky130_fd_sc_hd__dfxtp_1 _30212_ (.CLK(clknet_leaf_55_clk),
    .D(_00860_),
    .Q(\count_instr[51] ));
 sky130_fd_sc_hd__dfxtp_1 _30213_ (.CLK(clknet_leaf_55_clk),
    .D(_00861_),
    .Q(\count_instr[52] ));
 sky130_fd_sc_hd__dfxtp_1 _30214_ (.CLK(clknet_leaf_55_clk),
    .D(_00862_),
    .Q(\count_instr[53] ));
 sky130_fd_sc_hd__dfxtp_1 _30215_ (.CLK(clknet_leaf_54_clk),
    .D(_00863_),
    .Q(\count_instr[54] ));
 sky130_fd_sc_hd__dfxtp_1 _30216_ (.CLK(clknet_leaf_55_clk),
    .D(_00864_),
    .Q(\count_instr[55] ));
 sky130_fd_sc_hd__dfxtp_1 _30217_ (.CLK(clknet_leaf_55_clk),
    .D(_00865_),
    .Q(\count_instr[56] ));
 sky130_fd_sc_hd__dfxtp_1 _30218_ (.CLK(clknet_leaf_55_clk),
    .D(_00866_),
    .Q(\count_instr[57] ));
 sky130_fd_sc_hd__dfxtp_1 _30219_ (.CLK(clknet_leaf_55_clk),
    .D(_00867_),
    .Q(\count_instr[58] ));
 sky130_fd_sc_hd__dfxtp_1 _30220_ (.CLK(clknet_leaf_55_clk),
    .D(_00868_),
    .Q(\count_instr[59] ));
 sky130_fd_sc_hd__dfxtp_1 _30221_ (.CLK(clknet_leaf_57_clk),
    .D(_00869_),
    .Q(\count_instr[60] ));
 sky130_fd_sc_hd__dfxtp_1 _30222_ (.CLK(clknet_leaf_57_clk),
    .D(_00870_),
    .Q(\count_instr[61] ));
 sky130_fd_sc_hd__dfxtp_1 _30223_ (.CLK(clknet_leaf_57_clk),
    .D(_00871_),
    .Q(\count_instr[62] ));
 sky130_fd_sc_hd__dfxtp_1 _30224_ (.CLK(clknet_leaf_56_clk),
    .D(_00872_),
    .Q(\count_instr[63] ));
 sky130_fd_sc_hd__dfxtp_1 _30225_ (.CLK(clknet_leaf_91_clk),
    .D(_00873_),
    .Q(\reg_pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30226_ (.CLK(clknet_leaf_91_clk),
    .D(_00874_),
    .Q(\reg_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30227_ (.CLK(clknet_leaf_92_clk),
    .D(_00875_),
    .Q(\reg_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30228_ (.CLK(clknet_leaf_92_clk),
    .D(_00876_),
    .Q(\reg_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _30229_ (.CLK(clknet_leaf_92_clk),
    .D(_00877_),
    .Q(\reg_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _30230_ (.CLK(clknet_leaf_92_clk),
    .D(_00878_),
    .Q(\reg_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _30231_ (.CLK(clknet_leaf_92_clk),
    .D(_00879_),
    .Q(\reg_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _30232_ (.CLK(clknet_leaf_92_clk),
    .D(_00880_),
    .Q(\reg_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _30233_ (.CLK(clknet_leaf_25_clk),
    .D(_00881_),
    .Q(\reg_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _30234_ (.CLK(clknet_leaf_92_clk),
    .D(_00882_),
    .Q(\reg_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _30235_ (.CLK(clknet_leaf_22_clk),
    .D(_00883_),
    .Q(\reg_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _30236_ (.CLK(clknet_leaf_22_clk),
    .D(_00884_),
    .Q(\reg_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _30237_ (.CLK(clknet_leaf_22_clk),
    .D(_00885_),
    .Q(\reg_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _30238_ (.CLK(clknet_leaf_22_clk),
    .D(_00886_),
    .Q(\reg_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _30239_ (.CLK(clknet_leaf_22_clk),
    .D(_00887_),
    .Q(\reg_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _30240_ (.CLK(clknet_leaf_22_clk),
    .D(_00888_),
    .Q(\reg_pc[16] ));
 sky130_fd_sc_hd__dfxtp_1 _30241_ (.CLK(clknet_leaf_22_clk),
    .D(_00889_),
    .Q(\reg_pc[17] ));
 sky130_fd_sc_hd__dfxtp_1 _30242_ (.CLK(clknet_leaf_21_clk),
    .D(_00890_),
    .Q(\reg_pc[18] ));
 sky130_fd_sc_hd__dfxtp_1 _30243_ (.CLK(clknet_leaf_208_clk),
    .D(_00891_),
    .Q(\reg_pc[19] ));
 sky130_fd_sc_hd__dfxtp_1 _30244_ (.CLK(clknet_leaf_208_clk),
    .D(_00892_),
    .Q(\reg_pc[20] ));
 sky130_fd_sc_hd__dfxtp_1 _30245_ (.CLK(clknet_leaf_208_clk),
    .D(_00893_),
    .Q(\reg_pc[21] ));
 sky130_fd_sc_hd__dfxtp_1 _30246_ (.CLK(clknet_leaf_209_clk),
    .D(_00894_),
    .Q(\reg_pc[22] ));
 sky130_fd_sc_hd__dfxtp_1 _30247_ (.CLK(clknet_leaf_208_clk),
    .D(_00895_),
    .Q(\reg_pc[23] ));
 sky130_fd_sc_hd__dfxtp_1 _30248_ (.CLK(clknet_leaf_208_clk),
    .D(_00896_),
    .Q(\reg_pc[24] ));
 sky130_fd_sc_hd__dfxtp_1 _30249_ (.CLK(clknet_leaf_207_clk),
    .D(_00897_),
    .Q(\reg_pc[25] ));
 sky130_fd_sc_hd__dfxtp_1 _30250_ (.CLK(clknet_leaf_207_clk),
    .D(_00898_),
    .Q(\reg_pc[26] ));
 sky130_fd_sc_hd__dfxtp_1 _30251_ (.CLK(clknet_leaf_207_clk),
    .D(_00899_),
    .Q(\reg_pc[27] ));
 sky130_fd_sc_hd__dfxtp_2 _30252_ (.CLK(clknet_leaf_207_clk),
    .D(_00900_),
    .Q(\reg_pc[28] ));
 sky130_fd_sc_hd__dfxtp_1 _30253_ (.CLK(clknet_leaf_207_clk),
    .D(_00901_),
    .Q(\reg_pc[29] ));
 sky130_fd_sc_hd__dfxtp_1 _30254_ (.CLK(clknet_leaf_207_clk),
    .D(_00902_),
    .Q(\reg_pc[30] ));
 sky130_fd_sc_hd__dfxtp_2 _30255_ (.CLK(clknet_leaf_176_clk),
    .D(_00903_),
    .Q(\reg_pc[31] ));
 sky130_fd_sc_hd__dfxtp_1 _30256_ (.CLK(clknet_leaf_98_clk),
    .D(_00904_),
    .Q(\reg_next_pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30257_ (.CLK(clknet_leaf_95_clk),
    .D(_00905_),
    .Q(\reg_next_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30258_ (.CLK(clknet_leaf_95_clk),
    .D(_00906_),
    .Q(\reg_next_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30259_ (.CLK(clknet_leaf_94_clk),
    .D(_00907_),
    .Q(\reg_next_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _30260_ (.CLK(clknet_leaf_93_clk),
    .D(_00908_),
    .Q(\reg_next_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _30261_ (.CLK(clknet_leaf_93_clk),
    .D(_00909_),
    .Q(\reg_next_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _30262_ (.CLK(clknet_leaf_174_clk),
    .D(_00910_),
    .Q(\reg_next_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _30263_ (.CLK(clknet_leaf_93_clk),
    .D(_00911_),
    .Q(\reg_next_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _30264_ (.CLK(clknet_leaf_174_clk),
    .D(_00912_),
    .Q(\reg_next_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _30265_ (.CLK(clknet_leaf_174_clk),
    .D(_00913_),
    .Q(\reg_next_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _30266_ (.CLK(clknet_leaf_174_clk),
    .D(_00914_),
    .Q(\reg_next_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _30267_ (.CLK(clknet_leaf_174_clk),
    .D(_00915_),
    .Q(\reg_next_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _30268_ (.CLK(clknet_leaf_175_clk),
    .D(_00916_),
    .Q(\reg_next_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _30269_ (.CLK(clknet_leaf_174_clk),
    .D(_00917_),
    .Q(\reg_next_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _30270_ (.CLK(clknet_leaf_174_clk),
    .D(_00918_),
    .Q(\reg_next_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _30271_ (.CLK(clknet_leaf_175_clk),
    .D(_00919_),
    .Q(\reg_next_pc[16] ));
 sky130_fd_sc_hd__dfxtp_1 _30272_ (.CLK(clknet_leaf_176_clk),
    .D(_00920_),
    .Q(\reg_next_pc[17] ));
 sky130_fd_sc_hd__dfxtp_2 _30273_ (.CLK(clknet_leaf_205_clk),
    .D(_00921_),
    .Q(\reg_next_pc[18] ));
 sky130_fd_sc_hd__dfxtp_1 _30274_ (.CLK(clknet_leaf_205_clk),
    .D(_00922_),
    .Q(\reg_next_pc[19] ));
 sky130_fd_sc_hd__dfxtp_1 _30275_ (.CLK(clknet_leaf_201_clk),
    .D(_00923_),
    .Q(\reg_next_pc[20] ));
 sky130_fd_sc_hd__dfxtp_1 _30276_ (.CLK(clknet_leaf_201_clk),
    .D(_00924_),
    .Q(\reg_next_pc[21] ));
 sky130_fd_sc_hd__dfxtp_1 _30277_ (.CLK(clknet_leaf_205_clk),
    .D(_00925_),
    .Q(\reg_next_pc[22] ));
 sky130_fd_sc_hd__dfxtp_1 _30278_ (.CLK(clknet_leaf_205_clk),
    .D(_00926_),
    .Q(\reg_next_pc[23] ));
 sky130_fd_sc_hd__dfxtp_1 _30279_ (.CLK(clknet_5_17__leaf_clk),
    .D(_00927_),
    .Q(\reg_next_pc[24] ));
 sky130_fd_sc_hd__dfxtp_1 _30280_ (.CLK(clknet_leaf_201_clk),
    .D(_00928_),
    .Q(\reg_next_pc[25] ));
 sky130_fd_sc_hd__dfxtp_1 _30281_ (.CLK(clknet_5_17__leaf_clk),
    .D(_00929_),
    .Q(\reg_next_pc[26] ));
 sky130_fd_sc_hd__dfxtp_1 _30282_ (.CLK(clknet_leaf_177_clk),
    .D(_00930_),
    .Q(\reg_next_pc[27] ));
 sky130_fd_sc_hd__dfxtp_1 _30283_ (.CLK(clknet_leaf_177_clk),
    .D(_00931_),
    .Q(\reg_next_pc[28] ));
 sky130_fd_sc_hd__dfxtp_1 _30284_ (.CLK(clknet_leaf_177_clk),
    .D(_00932_),
    .Q(\reg_next_pc[29] ));
 sky130_fd_sc_hd__dfxtp_1 _30285_ (.CLK(clknet_leaf_177_clk),
    .D(_00933_),
    .Q(\reg_next_pc[30] ));
 sky130_fd_sc_hd__dfxtp_2 _30286_ (.CLK(clknet_leaf_172_clk),
    .D(_00934_),
    .Q(\reg_next_pc[31] ));
 sky130_fd_sc_hd__dfxtp_1 _30287_ (.CLK(clknet_leaf_67_clk),
    .D(_00935_),
    .Q(\count_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30288_ (.CLK(clknet_leaf_67_clk),
    .D(_00936_),
    .Q(\count_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30289_ (.CLK(clknet_leaf_67_clk),
    .D(_00937_),
    .Q(\count_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30290_ (.CLK(clknet_leaf_68_clk),
    .D(_00938_),
    .Q(\count_cycle[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30291_ (.CLK(clknet_leaf_68_clk),
    .D(_00939_),
    .Q(\count_cycle[4] ));
 sky130_fd_sc_hd__dfxtp_1 _30292_ (.CLK(clknet_leaf_68_clk),
    .D(_00940_),
    .Q(\count_cycle[5] ));
 sky130_fd_sc_hd__dfxtp_1 _30293_ (.CLK(clknet_leaf_68_clk),
    .D(_00941_),
    .Q(\count_cycle[6] ));
 sky130_fd_sc_hd__dfxtp_1 _30294_ (.CLK(clknet_leaf_65_clk),
    .D(_00942_),
    .Q(\count_cycle[7] ));
 sky130_fd_sc_hd__dfxtp_1 _30295_ (.CLK(clknet_leaf_65_clk),
    .D(_00943_),
    .Q(\count_cycle[8] ));
 sky130_fd_sc_hd__dfxtp_1 _30296_ (.CLK(clknet_leaf_66_clk),
    .D(_00944_),
    .Q(\count_cycle[9] ));
 sky130_fd_sc_hd__dfxtp_1 _30297_ (.CLK(clknet_leaf_63_clk),
    .D(_00945_),
    .Q(\count_cycle[10] ));
 sky130_fd_sc_hd__dfxtp_1 _30298_ (.CLK(clknet_leaf_63_clk),
    .D(_00946_),
    .Q(\count_cycle[11] ));
 sky130_fd_sc_hd__dfxtp_1 _30299_ (.CLK(clknet_leaf_63_clk),
    .D(_00947_),
    .Q(\count_cycle[12] ));
 sky130_fd_sc_hd__dfxtp_1 _30300_ (.CLK(clknet_leaf_63_clk),
    .D(_00948_),
    .Q(\count_cycle[13] ));
 sky130_fd_sc_hd__dfxtp_1 _30301_ (.CLK(clknet_leaf_63_clk),
    .D(_00949_),
    .Q(\count_cycle[14] ));
 sky130_fd_sc_hd__dfxtp_1 _30302_ (.CLK(clknet_leaf_63_clk),
    .D(_00950_),
    .Q(\count_cycle[15] ));
 sky130_fd_sc_hd__dfxtp_1 _30303_ (.CLK(clknet_leaf_50_clk),
    .D(_00951_),
    .Q(\count_cycle[16] ));
 sky130_fd_sc_hd__dfxtp_1 _30304_ (.CLK(clknet_leaf_63_clk),
    .D(_00952_),
    .Q(\count_cycle[17] ));
 sky130_fd_sc_hd__dfxtp_1 _30305_ (.CLK(clknet_leaf_51_clk),
    .D(_00953_),
    .Q(\count_cycle[18] ));
 sky130_fd_sc_hd__dfxtp_1 _30306_ (.CLK(clknet_leaf_51_clk),
    .D(_00954_),
    .Q(\count_cycle[19] ));
 sky130_fd_sc_hd__dfxtp_1 _30307_ (.CLK(clknet_leaf_51_clk),
    .D(_00955_),
    .Q(\count_cycle[20] ));
 sky130_fd_sc_hd__dfxtp_1 _30308_ (.CLK(clknet_leaf_51_clk),
    .D(_00956_),
    .Q(\count_cycle[21] ));
 sky130_fd_sc_hd__dfxtp_1 _30309_ (.CLK(clknet_leaf_62_clk),
    .D(_00957_),
    .Q(\count_cycle[22] ));
 sky130_fd_sc_hd__dfxtp_1 _30310_ (.CLK(clknet_leaf_63_clk),
    .D(_00958_),
    .Q(\count_cycle[23] ));
 sky130_fd_sc_hd__dfxtp_1 _30311_ (.CLK(clknet_leaf_62_clk),
    .D(_00959_),
    .Q(\count_cycle[24] ));
 sky130_fd_sc_hd__dfxtp_1 _30312_ (.CLK(clknet_leaf_61_clk),
    .D(_00960_),
    .Q(\count_cycle[25] ));
 sky130_fd_sc_hd__dfxtp_1 _30313_ (.CLK(clknet_leaf_60_clk),
    .D(_00961_),
    .Q(\count_cycle[26] ));
 sky130_fd_sc_hd__dfxtp_1 _30314_ (.CLK(clknet_leaf_60_clk),
    .D(_00962_),
    .Q(\count_cycle[27] ));
 sky130_fd_sc_hd__dfxtp_1 _30315_ (.CLK(clknet_leaf_59_clk),
    .D(_00963_),
    .Q(\count_cycle[28] ));
 sky130_fd_sc_hd__dfxtp_1 _30316_ (.CLK(clknet_leaf_59_clk),
    .D(_00964_),
    .Q(\count_cycle[29] ));
 sky130_fd_sc_hd__dfxtp_1 _30317_ (.CLK(clknet_leaf_59_clk),
    .D(_00965_),
    .Q(\count_cycle[30] ));
 sky130_fd_sc_hd__dfxtp_1 _30318_ (.CLK(clknet_leaf_70_clk),
    .D(_00966_),
    .Q(\count_cycle[31] ));
 sky130_fd_sc_hd__dfxtp_1 _30319_ (.CLK(clknet_leaf_70_clk),
    .D(_00967_),
    .Q(\count_cycle[32] ));
 sky130_fd_sc_hd__dfxtp_1 _30320_ (.CLK(clknet_leaf_70_clk),
    .D(_00968_),
    .Q(\count_cycle[33] ));
 sky130_fd_sc_hd__dfxtp_1 _30321_ (.CLK(clknet_leaf_70_clk),
    .D(_00969_),
    .Q(\count_cycle[34] ));
 sky130_fd_sc_hd__dfxtp_1 _30322_ (.CLK(clknet_leaf_71_clk),
    .D(_00970_),
    .Q(\count_cycle[35] ));
 sky130_fd_sc_hd__dfxtp_1 _30323_ (.CLK(clknet_leaf_70_clk),
    .D(_00971_),
    .Q(\count_cycle[36] ));
 sky130_fd_sc_hd__dfxtp_1 _30324_ (.CLK(clknet_leaf_69_clk),
    .D(_00972_),
    .Q(\count_cycle[37] ));
 sky130_fd_sc_hd__dfxtp_1 _30325_ (.CLK(clknet_leaf_69_clk),
    .D(_00973_),
    .Q(\count_cycle[38] ));
 sky130_fd_sc_hd__dfxtp_1 _30326_ (.CLK(clknet_leaf_69_clk),
    .D(_00974_),
    .Q(\count_cycle[39] ));
 sky130_fd_sc_hd__dfxtp_1 _30327_ (.CLK(clknet_leaf_69_clk),
    .D(_00975_),
    .Q(\count_cycle[40] ));
 sky130_fd_sc_hd__dfxtp_1 _30328_ (.CLK(clknet_leaf_69_clk),
    .D(_00976_),
    .Q(\count_cycle[41] ));
 sky130_fd_sc_hd__dfxtp_1 _30329_ (.CLK(clknet_leaf_59_clk),
    .D(_00977_),
    .Q(\count_cycle[42] ));
 sky130_fd_sc_hd__dfxtp_1 _30330_ (.CLK(clknet_leaf_59_clk),
    .D(_00978_),
    .Q(\count_cycle[43] ));
 sky130_fd_sc_hd__dfxtp_1 _30331_ (.CLK(clknet_leaf_59_clk),
    .D(_00979_),
    .Q(\count_cycle[44] ));
 sky130_fd_sc_hd__dfxtp_1 _30332_ (.CLK(clknet_leaf_58_clk),
    .D(_00980_),
    .Q(\count_cycle[45] ));
 sky130_fd_sc_hd__dfxtp_1 _30333_ (.CLK(clknet_leaf_58_clk),
    .D(_00981_),
    .Q(\count_cycle[46] ));
 sky130_fd_sc_hd__dfxtp_1 _30334_ (.CLK(clknet_leaf_57_clk),
    .D(_00982_),
    .Q(\count_cycle[47] ));
 sky130_fd_sc_hd__dfxtp_1 _30335_ (.CLK(clknet_leaf_56_clk),
    .D(_00983_),
    .Q(\count_cycle[48] ));
 sky130_fd_sc_hd__dfxtp_1 _30336_ (.CLK(clknet_leaf_56_clk),
    .D(_00984_),
    .Q(\count_cycle[49] ));
 sky130_fd_sc_hd__dfxtp_1 _30337_ (.CLK(clknet_leaf_54_clk),
    .D(_00985_),
    .Q(\count_cycle[50] ));
 sky130_fd_sc_hd__dfxtp_1 _30338_ (.CLK(clknet_leaf_54_clk),
    .D(_00986_),
    .Q(\count_cycle[51] ));
 sky130_fd_sc_hd__dfxtp_1 _30339_ (.CLK(clknet_leaf_54_clk),
    .D(_00987_),
    .Q(\count_cycle[52] ));
 sky130_fd_sc_hd__dfxtp_1 _30340_ (.CLK(clknet_leaf_54_clk),
    .D(_00988_),
    .Q(\count_cycle[53] ));
 sky130_fd_sc_hd__dfxtp_1 _30341_ (.CLK(clknet_leaf_54_clk),
    .D(_00989_),
    .Q(\count_cycle[54] ));
 sky130_fd_sc_hd__dfxtp_1 _30342_ (.CLK(clknet_leaf_52_clk),
    .D(_00990_),
    .Q(\count_cycle[55] ));
 sky130_fd_sc_hd__dfxtp_1 _30343_ (.CLK(clknet_leaf_54_clk),
    .D(_00991_),
    .Q(\count_cycle[56] ));
 sky130_fd_sc_hd__dfxtp_1 _30344_ (.CLK(clknet_leaf_52_clk),
    .D(_00992_),
    .Q(\count_cycle[57] ));
 sky130_fd_sc_hd__dfxtp_1 _30345_ (.CLK(clknet_leaf_52_clk),
    .D(_00993_),
    .Q(\count_cycle[58] ));
 sky130_fd_sc_hd__dfxtp_1 _30346_ (.CLK(clknet_leaf_54_clk),
    .D(_00994_),
    .Q(\count_cycle[59] ));
 sky130_fd_sc_hd__dfxtp_1 _30347_ (.CLK(clknet_leaf_62_clk),
    .D(_00995_),
    .Q(\count_cycle[60] ));
 sky130_fd_sc_hd__dfxtp_1 _30348_ (.CLK(clknet_leaf_51_clk),
    .D(_00996_),
    .Q(\count_cycle[61] ));
 sky130_fd_sc_hd__dfxtp_1 _30349_ (.CLK(clknet_leaf_51_clk),
    .D(_00997_),
    .Q(\count_cycle[62] ));
 sky130_fd_sc_hd__dfxtp_1 _30350_ (.CLK(clknet_leaf_51_clk),
    .D(_00998_),
    .Q(\count_cycle[63] ));
 sky130_fd_sc_hd__dfxtp_2 _30351_ (.CLK(clknet_leaf_33_clk),
    .D(_00999_),
    .Q(net267));
 sky130_fd_sc_hd__dfxtp_4 _30352_ (.CLK(clknet_leaf_33_clk),
    .D(_01000_),
    .Q(net278));
 sky130_fd_sc_hd__dfxtp_1 _30353_ (.CLK(clknet_leaf_33_clk),
    .D(_01001_),
    .Q(net289));
 sky130_fd_sc_hd__dfxtp_2 _30354_ (.CLK(clknet_leaf_34_clk),
    .D(_01002_),
    .Q(net292));
 sky130_fd_sc_hd__dfxtp_4 _30355_ (.CLK(clknet_leaf_28_clk),
    .D(_01003_),
    .Q(net293));
 sky130_fd_sc_hd__dfxtp_2 _30356_ (.CLK(clknet_leaf_35_clk),
    .D(_01004_),
    .Q(net294));
 sky130_fd_sc_hd__dfxtp_2 _30357_ (.CLK(clknet_leaf_35_clk),
    .D(_01005_),
    .Q(net295));
 sky130_fd_sc_hd__dfxtp_2 _30358_ (.CLK(clknet_leaf_35_clk),
    .D(_01006_),
    .Q(net296));
 sky130_fd_sc_hd__dfxtp_2 _30359_ (.CLK(clknet_leaf_35_clk),
    .D(_01007_),
    .Q(net297));
 sky130_fd_sc_hd__dfxtp_2 _30360_ (.CLK(clknet_leaf_36_clk),
    .D(_01008_),
    .Q(net298));
 sky130_fd_sc_hd__dfxtp_2 _30361_ (.CLK(clknet_leaf_27_clk),
    .D(_01009_),
    .Q(net268));
 sky130_fd_sc_hd__dfxtp_2 _30362_ (.CLK(clknet_leaf_20_clk),
    .D(_01010_),
    .Q(net269));
 sky130_fd_sc_hd__dfxtp_2 _30363_ (.CLK(clknet_leaf_20_clk),
    .D(_01011_),
    .Q(net270));
 sky130_fd_sc_hd__dfxtp_2 _30364_ (.CLK(clknet_leaf_20_clk),
    .D(_01012_),
    .Q(net271));
 sky130_fd_sc_hd__dfxtp_2 _30365_ (.CLK(clknet_leaf_20_clk),
    .D(_01013_),
    .Q(net272));
 sky130_fd_sc_hd__dfxtp_4 _30366_ (.CLK(clknet_leaf_19_clk),
    .D(_01014_),
    .Q(net273));
 sky130_fd_sc_hd__dfxtp_4 _30367_ (.CLK(clknet_leaf_19_clk),
    .D(_01015_),
    .Q(net274));
 sky130_fd_sc_hd__dfxtp_2 _30368_ (.CLK(clknet_leaf_19_clk),
    .D(_01016_),
    .Q(net275));
 sky130_fd_sc_hd__dfxtp_4 _30369_ (.CLK(clknet_leaf_19_clk),
    .D(_01017_),
    .Q(net276));
 sky130_fd_sc_hd__dfxtp_2 _30370_ (.CLK(clknet_leaf_18_clk),
    .D(_01018_),
    .Q(net277));
 sky130_fd_sc_hd__dfxtp_4 _30371_ (.CLK(clknet_leaf_17_clk),
    .D(_01019_),
    .Q(net279));
 sky130_fd_sc_hd__dfxtp_4 _30372_ (.CLK(clknet_leaf_17_clk),
    .D(_01020_),
    .Q(net280));
 sky130_fd_sc_hd__dfxtp_4 _30373_ (.CLK(clknet_leaf_17_clk),
    .D(_01021_),
    .Q(net281));
 sky130_fd_sc_hd__dfxtp_2 _30374_ (.CLK(clknet_leaf_17_clk),
    .D(_01022_),
    .Q(net282));
 sky130_fd_sc_hd__dfxtp_2 _30375_ (.CLK(clknet_leaf_15_clk),
    .D(_01023_),
    .Q(net283));
 sky130_fd_sc_hd__dfxtp_2 _30376_ (.CLK(clknet_leaf_15_clk),
    .D(_01024_),
    .Q(net284));
 sky130_fd_sc_hd__dfxtp_2 _30377_ (.CLK(clknet_leaf_15_clk),
    .D(_01025_),
    .Q(net285));
 sky130_fd_sc_hd__dfxtp_4 _30378_ (.CLK(clknet_leaf_13_clk),
    .D(_01026_),
    .Q(net286));
 sky130_fd_sc_hd__dfxtp_2 _30379_ (.CLK(clknet_leaf_19_clk),
    .D(_01027_),
    .Q(net287));
 sky130_fd_sc_hd__dfxtp_4 _30380_ (.CLK(clknet_leaf_19_clk),
    .D(_01028_),
    .Q(net288));
 sky130_fd_sc_hd__dfxtp_2 _30381_ (.CLK(clknet_leaf_19_clk),
    .D(_01029_),
    .Q(net290));
 sky130_fd_sc_hd__dfxtp_2 _30382_ (.CLK(clknet_leaf_13_clk),
    .D(_01030_),
    .Q(net291));
 sky130_fd_sc_hd__dfxtp_1 _30383_ (.CLK(clknet_leaf_82_clk),
    .D(_14572_),
    .Q(\reg_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30384_ (.CLK(clknet_leaf_83_clk),
    .D(_14583_),
    .Q(\reg_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30385_ (.CLK(clknet_leaf_82_clk),
    .D(_14594_),
    .Q(\reg_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30386_ (.CLK(clknet_leaf_79_clk),
    .D(_14597_),
    .Q(\reg_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30387_ (.CLK(clknet_leaf_91_clk),
    .D(_14598_),
    .Q(\reg_out[4] ));
 sky130_fd_sc_hd__dfxtp_1 _30388_ (.CLK(clknet_leaf_82_clk),
    .D(_14599_),
    .Q(\reg_out[5] ));
 sky130_fd_sc_hd__dfxtp_1 _30389_ (.CLK(clknet_leaf_89_clk),
    .D(_14600_),
    .Q(\reg_out[6] ));
 sky130_fd_sc_hd__dfxtp_1 _30390_ (.CLK(clknet_leaf_92_clk),
    .D(_14601_),
    .Q(\reg_out[7] ));
 sky130_fd_sc_hd__dfxtp_1 _30391_ (.CLK(clknet_leaf_23_clk),
    .D(_14602_),
    .Q(\reg_out[8] ));
 sky130_fd_sc_hd__dfxtp_1 _30392_ (.CLK(clknet_leaf_23_clk),
    .D(_14603_),
    .Q(\reg_out[9] ));
 sky130_fd_sc_hd__dfxtp_1 _30393_ (.CLK(clknet_leaf_23_clk),
    .D(_14573_),
    .Q(\reg_out[10] ));
 sky130_fd_sc_hd__dfxtp_1 _30394_ (.CLK(clknet_leaf_23_clk),
    .D(_14574_),
    .Q(\reg_out[11] ));
 sky130_fd_sc_hd__dfxtp_1 _30395_ (.CLK(clknet_leaf_23_clk),
    .D(_14575_),
    .Q(\reg_out[12] ));
 sky130_fd_sc_hd__dfxtp_1 _30396_ (.CLK(clknet_leaf_23_clk),
    .D(_14576_),
    .Q(\reg_out[13] ));
 sky130_fd_sc_hd__dfxtp_1 _30397_ (.CLK(clknet_leaf_23_clk),
    .D(_14577_),
    .Q(\reg_out[14] ));
 sky130_fd_sc_hd__dfxtp_1 _30398_ (.CLK(clknet_leaf_23_clk),
    .D(_14578_),
    .Q(\reg_out[15] ));
 sky130_fd_sc_hd__dfxtp_1 _30399_ (.CLK(clknet_leaf_21_clk),
    .D(_14579_),
    .Q(\reg_out[16] ));
 sky130_fd_sc_hd__dfxtp_1 _30400_ (.CLK(clknet_leaf_23_clk),
    .D(_14580_),
    .Q(\reg_out[17] ));
 sky130_fd_sc_hd__dfxtp_1 _30401_ (.CLK(clknet_leaf_209_clk),
    .D(_14581_),
    .Q(\reg_out[18] ));
 sky130_fd_sc_hd__dfxtp_1 _30402_ (.CLK(clknet_leaf_209_clk),
    .D(_14582_),
    .Q(\reg_out[19] ));
 sky130_fd_sc_hd__dfxtp_1 _30403_ (.CLK(clknet_leaf_209_clk),
    .D(_14584_),
    .Q(\reg_out[20] ));
 sky130_fd_sc_hd__dfxtp_1 _30404_ (.CLK(clknet_leaf_209_clk),
    .D(_14585_),
    .Q(\reg_out[21] ));
 sky130_fd_sc_hd__dfxtp_1 _30405_ (.CLK(clknet_leaf_209_clk),
    .D(_14586_),
    .Q(\reg_out[22] ));
 sky130_fd_sc_hd__dfxtp_1 _30406_ (.CLK(clknet_leaf_209_clk),
    .D(_14587_),
    .Q(\reg_out[23] ));
 sky130_fd_sc_hd__dfxtp_1 _30407_ (.CLK(clknet_leaf_209_clk),
    .D(_14588_),
    .Q(\reg_out[24] ));
 sky130_fd_sc_hd__dfxtp_1 _30408_ (.CLK(clknet_leaf_208_clk),
    .D(_14589_),
    .Q(\reg_out[25] ));
 sky130_fd_sc_hd__dfxtp_1 _30409_ (.CLK(clknet_leaf_209_clk),
    .D(_14590_),
    .Q(\reg_out[26] ));
 sky130_fd_sc_hd__dfxtp_1 _30410_ (.CLK(clknet_leaf_21_clk),
    .D(_14591_),
    .Q(\reg_out[27] ));
 sky130_fd_sc_hd__dfxtp_1 _30411_ (.CLK(clknet_leaf_21_clk),
    .D(_14592_),
    .Q(\reg_out[28] ));
 sky130_fd_sc_hd__dfxtp_1 _30412_ (.CLK(clknet_leaf_21_clk),
    .D(_14593_),
    .Q(\reg_out[29] ));
 sky130_fd_sc_hd__dfxtp_1 _30413_ (.CLK(clknet_leaf_21_clk),
    .D(_14595_),
    .Q(\reg_out[30] ));
 sky130_fd_sc_hd__dfxtp_1 _30414_ (.CLK(clknet_leaf_21_clk),
    .D(_14596_),
    .Q(\reg_out[31] ));
 sky130_fd_sc_hd__dfxtp_1 _30415_ (.CLK(clknet_leaf_81_clk),
    .D(_01031_),
    .Q(irq_delay));
 sky130_fd_sc_hd__dfxtp_1 _30416_ (.CLK(clknet_leaf_81_clk),
    .D(_01032_),
    .Q(irq_active));
 sky130_fd_sc_hd__dfxtp_1 _30417_ (.CLK(clknet_leaf_74_clk),
    .D(_01033_),
    .Q(\irq_mask[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30418_ (.CLK(clknet_leaf_74_clk),
    .D(_01034_),
    .Q(\irq_mask[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30419_ (.CLK(clknet_leaf_74_clk),
    .D(_01035_),
    .Q(\irq_mask[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30420_ (.CLK(clknet_leaf_74_clk),
    .D(_01036_),
    .Q(\irq_mask[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30421_ (.CLK(clknet_leaf_75_clk),
    .D(_01037_),
    .Q(\irq_mask[4] ));
 sky130_fd_sc_hd__dfxtp_1 _30422_ (.CLK(clknet_leaf_73_clk),
    .D(_01038_),
    .Q(\irq_mask[5] ));
 sky130_fd_sc_hd__dfxtp_1 _30423_ (.CLK(clknet_leaf_77_clk),
    .D(_01039_),
    .Q(\irq_mask[6] ));
 sky130_fd_sc_hd__dfxtp_1 _30424_ (.CLK(clknet_leaf_78_clk),
    .D(_01040_),
    .Q(\irq_mask[7] ));
 sky130_fd_sc_hd__dfxtp_1 _30425_ (.CLK(clknet_leaf_78_clk),
    .D(_01041_),
    .Q(\irq_mask[8] ));
 sky130_fd_sc_hd__dfxtp_1 _30426_ (.CLK(clknet_leaf_77_clk),
    .D(_01042_),
    .Q(\irq_mask[9] ));
 sky130_fd_sc_hd__dfxtp_1 _30427_ (.CLK(clknet_leaf_78_clk),
    .D(_01043_),
    .Q(\irq_mask[10] ));
 sky130_fd_sc_hd__dfxtp_1 _30428_ (.CLK(clknet_leaf_79_clk),
    .D(_01044_),
    .Q(\irq_mask[11] ));
 sky130_fd_sc_hd__dfxtp_1 _30429_ (.CLK(clknet_leaf_79_clk),
    .D(_01045_),
    .Q(\irq_mask[12] ));
 sky130_fd_sc_hd__dfxtp_1 _30430_ (.CLK(clknet_leaf_80_clk),
    .D(_01046_),
    .Q(\irq_mask[13] ));
 sky130_fd_sc_hd__dfxtp_1 _30431_ (.CLK(clknet_leaf_80_clk),
    .D(_01047_),
    .Q(\irq_mask[14] ));
 sky130_fd_sc_hd__dfxtp_1 _30432_ (.CLK(clknet_leaf_111_clk),
    .D(_01048_),
    .Q(\irq_mask[15] ));
 sky130_fd_sc_hd__dfxtp_1 _30433_ (.CLK(clknet_leaf_111_clk),
    .D(_01049_),
    .Q(\irq_mask[16] ));
 sky130_fd_sc_hd__dfxtp_1 _30434_ (.CLK(clknet_leaf_108_clk),
    .D(_01050_),
    .Q(\irq_mask[17] ));
 sky130_fd_sc_hd__dfxtp_1 _30435_ (.CLK(clknet_leaf_111_clk),
    .D(_01051_),
    .Q(\irq_mask[18] ));
 sky130_fd_sc_hd__dfxtp_1 _30436_ (.CLK(clknet_leaf_77_clk),
    .D(_01052_),
    .Q(\irq_mask[19] ));
 sky130_fd_sc_hd__dfxtp_1 _30437_ (.CLK(clknet_leaf_112_clk),
    .D(_01053_),
    .Q(\irq_mask[20] ));
 sky130_fd_sc_hd__dfxtp_1 _30438_ (.CLK(clknet_leaf_111_clk),
    .D(_01054_),
    .Q(\irq_mask[21] ));
 sky130_fd_sc_hd__dfxtp_1 _30439_ (.CLK(clknet_leaf_76_clk),
    .D(_01055_),
    .Q(\irq_mask[22] ));
 sky130_fd_sc_hd__dfxtp_1 _30440_ (.CLK(clknet_leaf_112_clk),
    .D(_01056_),
    .Q(\irq_mask[23] ));
 sky130_fd_sc_hd__dfxtp_1 _30441_ (.CLK(clknet_leaf_76_clk),
    .D(_01057_),
    .Q(\irq_mask[24] ));
 sky130_fd_sc_hd__dfxtp_2 _30442_ (.CLK(clknet_leaf_75_clk),
    .D(_01058_),
    .Q(\irq_mask[25] ));
 sky130_fd_sc_hd__dfxtp_1 _30443_ (.CLK(clknet_leaf_76_clk),
    .D(_01059_),
    .Q(\irq_mask[26] ));
 sky130_fd_sc_hd__dfxtp_1 _30444_ (.CLK(clknet_leaf_75_clk),
    .D(_01060_),
    .Q(\irq_mask[27] ));
 sky130_fd_sc_hd__dfxtp_1 _30445_ (.CLK(clknet_leaf_75_clk),
    .D(_01061_),
    .Q(\irq_mask[28] ));
 sky130_fd_sc_hd__dfxtp_1 _30446_ (.CLK(clknet_leaf_75_clk),
    .D(_01062_),
    .Q(\irq_mask[29] ));
 sky130_fd_sc_hd__dfxtp_1 _30447_ (.CLK(clknet_leaf_75_clk),
    .D(_01063_),
    .Q(\irq_mask[30] ));
 sky130_fd_sc_hd__dfxtp_1 _30448_ (.CLK(clknet_leaf_73_clk),
    .D(_01064_),
    .Q(\irq_mask[31] ));
 sky130_fd_sc_hd__dfxtp_4 _30449_ (.CLK(clknet_leaf_35_clk),
    .D(_01065_),
    .Q(net161));
 sky130_fd_sc_hd__dfxtp_2 _30450_ (.CLK(clknet_leaf_34_clk),
    .D(_01066_),
    .Q(net172));
 sky130_fd_sc_hd__dfxtp_1 _30451_ (.CLK(clknet_leaf_34_clk),
    .D(_01067_),
    .Q(net183));
 sky130_fd_sc_hd__dfxtp_2 _30452_ (.CLK(clknet_leaf_34_clk),
    .D(_01068_),
    .Q(net186));
 sky130_fd_sc_hd__dfxtp_2 _30453_ (.CLK(clknet_leaf_34_clk),
    .D(_01069_),
    .Q(net187));
 sky130_fd_sc_hd__dfxtp_2 _30454_ (.CLK(clknet_leaf_35_clk),
    .D(_01070_),
    .Q(net188));
 sky130_fd_sc_hd__dfxtp_2 _30455_ (.CLK(clknet_leaf_35_clk),
    .D(_01071_),
    .Q(net189));
 sky130_fd_sc_hd__dfxtp_2 _30456_ (.CLK(clknet_leaf_35_clk),
    .D(_01072_),
    .Q(net190));
 sky130_fd_sc_hd__dfxtp_1 _30457_ (.CLK(clknet_leaf_36_clk),
    .D(_01073_),
    .Q(net329));
 sky130_fd_sc_hd__dfxtp_2 _30458_ (.CLK(clknet_leaf_36_clk),
    .D(_01074_),
    .Q(net330));
 sky130_fd_sc_hd__dfxtp_1 _30459_ (.CLK(clknet_leaf_36_clk),
    .D(_01075_),
    .Q(net300));
 sky130_fd_sc_hd__dfxtp_2 _30460_ (.CLK(clknet_leaf_12_clk),
    .D(_01076_),
    .Q(net301));
 sky130_fd_sc_hd__dfxtp_4 _30461_ (.CLK(clknet_leaf_12_clk),
    .D(_01077_),
    .Q(net302));
 sky130_fd_sc_hd__dfxtp_2 _30462_ (.CLK(clknet_leaf_12_clk),
    .D(_01078_),
    .Q(net303));
 sky130_fd_sc_hd__dfxtp_2 _30463_ (.CLK(clknet_leaf_12_clk),
    .D(_01079_),
    .Q(net304));
 sky130_fd_sc_hd__dfxtp_2 _30464_ (.CLK(clknet_leaf_12_clk),
    .D(_01080_),
    .Q(net305));
 sky130_fd_sc_hd__dfxtp_4 _30465_ (.CLK(clknet_leaf_12_clk),
    .D(_01081_),
    .Q(net306));
 sky130_fd_sc_hd__dfxtp_2 _30466_ (.CLK(clknet_leaf_15_clk),
    .D(_01082_),
    .Q(net307));
 sky130_fd_sc_hd__dfxtp_4 _30467_ (.CLK(clknet_leaf_13_clk),
    .D(_01083_),
    .Q(net308));
 sky130_fd_sc_hd__dfxtp_2 _30468_ (.CLK(clknet_leaf_15_clk),
    .D(_01084_),
    .Q(net309));
 sky130_fd_sc_hd__dfxtp_2 _30469_ (.CLK(clknet_leaf_16_clk),
    .D(_01085_),
    .Q(net311));
 sky130_fd_sc_hd__dfxtp_2 _30470_ (.CLK(clknet_leaf_16_clk),
    .D(_01086_),
    .Q(net312));
 sky130_fd_sc_hd__dfxtp_4 _30471_ (.CLK(clknet_leaf_15_clk),
    .D(_01087_),
    .Q(net313));
 sky130_fd_sc_hd__dfxtp_2 _30472_ (.CLK(clknet_leaf_15_clk),
    .D(_01088_),
    .Q(net314));
 sky130_fd_sc_hd__dfxtp_4 _30473_ (.CLK(clknet_leaf_13_clk),
    .D(_01089_),
    .Q(net315));
 sky130_fd_sc_hd__dfxtp_1 _30474_ (.CLK(clknet_leaf_15_clk),
    .D(_01090_),
    .Q(net316));
 sky130_fd_sc_hd__dfxtp_4 _30475_ (.CLK(clknet_leaf_19_clk),
    .D(_01091_),
    .Q(net317));
 sky130_fd_sc_hd__dfxtp_2 _30476_ (.CLK(clknet_leaf_13_clk),
    .D(_01092_),
    .Q(net318));
 sky130_fd_sc_hd__dfxtp_2 _30477_ (.CLK(clknet_leaf_13_clk),
    .D(_01093_),
    .Q(net319));
 sky130_fd_sc_hd__dfxtp_4 _30478_ (.CLK(clknet_leaf_13_clk),
    .D(_01094_),
    .Q(net320));
 sky130_fd_sc_hd__dfxtp_2 _30479_ (.CLK(clknet_leaf_13_clk),
    .D(_01095_),
    .Q(net322));
 sky130_fd_sc_hd__dfxtp_2 _30480_ (.CLK(clknet_leaf_12_clk),
    .D(_01096_),
    .Q(net323));
 sky130_fd_sc_hd__dfxtp_1 _30481_ (.CLK(clknet_leaf_79_clk),
    .D(_01097_),
    .Q(\irq_pending[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30482_ (.CLK(clknet_leaf_83_clk),
    .D(_01098_),
    .Q(\irq_pending[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30483_ (.CLK(clknet_leaf_79_clk),
    .D(_01099_),
    .Q(\irq_pending[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30484_ (.CLK(clknet_leaf_79_clk),
    .D(_01100_),
    .Q(\irq_pending[4] ));
 sky130_fd_sc_hd__dfxtp_1 _30485_ (.CLK(clknet_leaf_79_clk),
    .D(_01101_),
    .Q(\irq_pending[5] ));
 sky130_fd_sc_hd__dfxtp_1 _30486_ (.CLK(clknet_leaf_79_clk),
    .D(_01102_),
    .Q(\irq_pending[6] ));
 sky130_fd_sc_hd__dfxtp_1 _30487_ (.CLK(clknet_leaf_79_clk),
    .D(_01103_),
    .Q(\irq_pending[7] ));
 sky130_fd_sc_hd__dfxtp_1 _30488_ (.CLK(clknet_leaf_80_clk),
    .D(_01104_),
    .Q(\irq_pending[8] ));
 sky130_fd_sc_hd__dfxtp_1 _30489_ (.CLK(clknet_leaf_80_clk),
    .D(_01105_),
    .Q(\irq_pending[9] ));
 sky130_fd_sc_hd__dfxtp_1 _30490_ (.CLK(clknet_leaf_80_clk),
    .D(_01106_),
    .Q(\irq_pending[10] ));
 sky130_fd_sc_hd__dfxtp_1 _30491_ (.CLK(clknet_leaf_80_clk),
    .D(_01107_),
    .Q(\irq_pending[11] ));
 sky130_fd_sc_hd__dfxtp_1 _30492_ (.CLK(clknet_leaf_80_clk),
    .D(_01108_),
    .Q(\irq_pending[12] ));
 sky130_fd_sc_hd__dfxtp_1 _30493_ (.CLK(clknet_leaf_80_clk),
    .D(_01109_),
    .Q(\irq_pending[13] ));
 sky130_fd_sc_hd__dfxtp_1 _30494_ (.CLK(clknet_leaf_90_clk),
    .D(_01110_),
    .Q(\irq_pending[14] ));
 sky130_fd_sc_hd__dfxtp_1 _30495_ (.CLK(clknet_leaf_90_clk),
    .D(_01111_),
    .Q(\irq_pending[15] ));
 sky130_fd_sc_hd__dfxtp_1 _30496_ (.CLK(clknet_leaf_81_clk),
    .D(_01112_),
    .Q(\irq_pending[16] ));
 sky130_fd_sc_hd__dfxtp_1 _30497_ (.CLK(clknet_leaf_90_clk),
    .D(_01113_),
    .Q(\irq_pending[17] ));
 sky130_fd_sc_hd__dfxtp_1 _30498_ (.CLK(clknet_leaf_90_clk),
    .D(_01114_),
    .Q(\irq_pending[18] ));
 sky130_fd_sc_hd__dfxtp_1 _30499_ (.CLK(clknet_leaf_90_clk),
    .D(_01115_),
    .Q(\irq_pending[19] ));
 sky130_fd_sc_hd__dfxtp_1 _30500_ (.CLK(clknet_leaf_95_clk),
    .D(_01116_),
    .Q(\irq_pending[20] ));
 sky130_fd_sc_hd__dfxtp_1 _30501_ (.CLK(clknet_leaf_96_clk),
    .D(_01117_),
    .Q(\irq_pending[21] ));
 sky130_fd_sc_hd__dfxtp_1 _30502_ (.CLK(clknet_leaf_95_clk),
    .D(_01118_),
    .Q(\irq_pending[22] ));
 sky130_fd_sc_hd__dfxtp_1 _30503_ (.CLK(clknet_leaf_107_clk),
    .D(_01119_),
    .Q(\irq_pending[23] ));
 sky130_fd_sc_hd__dfxtp_1 _30504_ (.CLK(clknet_leaf_107_clk),
    .D(_01120_),
    .Q(\irq_pending[24] ));
 sky130_fd_sc_hd__dfxtp_1 _30505_ (.CLK(clknet_leaf_81_clk),
    .D(_01121_),
    .Q(\irq_pending[25] ));
 sky130_fd_sc_hd__dfxtp_1 _30506_ (.CLK(clknet_leaf_107_clk),
    .D(_01122_),
    .Q(\irq_pending[26] ));
 sky130_fd_sc_hd__dfxtp_1 _30507_ (.CLK(clknet_leaf_107_clk),
    .D(_01123_),
    .Q(\irq_pending[27] ));
 sky130_fd_sc_hd__dfxtp_1 _30508_ (.CLK(clknet_leaf_80_clk),
    .D(_01124_),
    .Q(\irq_pending[28] ));
 sky130_fd_sc_hd__dfxtp_1 _30509_ (.CLK(clknet_leaf_80_clk),
    .D(_01125_),
    .Q(\irq_pending[29] ));
 sky130_fd_sc_hd__dfxtp_1 _30510_ (.CLK(clknet_leaf_108_clk),
    .D(_01126_),
    .Q(\irq_pending[30] ));
 sky130_fd_sc_hd__dfxtp_1 _30511_ (.CLK(clknet_leaf_80_clk),
    .D(_01127_),
    .Q(\irq_pending[31] ));
 sky130_fd_sc_hd__dfxtp_1 _30512_ (.CLK(clknet_leaf_85_clk),
    .D(_01128_),
    .Q(mem_do_prefetch));
 sky130_fd_sc_hd__dfxtp_1 _30513_ (.CLK(clknet_leaf_89_clk),
    .D(_01129_),
    .Q(mem_do_rinst));
 sky130_fd_sc_hd__dfxtp_1 _30514_ (.CLK(clknet_leaf_84_clk),
    .D(_01130_),
    .Q(mem_do_rdata));
 sky130_fd_sc_hd__dfxtp_1 _30515_ (.CLK(clknet_leaf_82_clk),
    .D(_01131_),
    .Q(mem_do_wdata));
 sky130_fd_sc_hd__dfxtp_1 _30516_ (.CLK(clknet_leaf_96_clk),
    .D(_00035_),
    .Q(decoder_trigger));
 sky130_fd_sc_hd__dfxtp_1 _30517_ (.CLK(clknet_leaf_112_clk),
    .D(_01132_),
    .Q(\timer[0] ));
 sky130_fd_sc_hd__dfxtp_2 _30518_ (.CLK(clknet_leaf_113_clk),
    .D(_01133_),
    .Q(\timer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30519_ (.CLK(clknet_leaf_112_clk),
    .D(_01134_),
    .Q(\timer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30520_ (.CLK(clknet_leaf_111_clk),
    .D(_01135_),
    .Q(\timer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30521_ (.CLK(clknet_leaf_111_clk),
    .D(_01136_),
    .Q(\timer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _30522_ (.CLK(clknet_leaf_108_clk),
    .D(_01137_),
    .Q(\timer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _30523_ (.CLK(clknet_leaf_108_clk),
    .D(_01138_),
    .Q(\timer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _30524_ (.CLK(clknet_leaf_109_clk),
    .D(_01139_),
    .Q(\timer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _30525_ (.CLK(clknet_leaf_110_clk),
    .D(_01140_),
    .Q(\timer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _30526_ (.CLK(clknet_leaf_111_clk),
    .D(_01141_),
    .Q(\timer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _30527_ (.CLK(clknet_leaf_114_clk),
    .D(_01142_),
    .Q(\timer[10] ));
 sky130_fd_sc_hd__dfxtp_2 _30528_ (.CLK(clknet_leaf_114_clk),
    .D(_01143_),
    .Q(\timer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _30529_ (.CLK(clknet_leaf_110_clk),
    .D(_01144_),
    .Q(\timer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _30530_ (.CLK(clknet_leaf_109_clk),
    .D(_01145_),
    .Q(\timer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _30531_ (.CLK(clknet_leaf_109_clk),
    .D(_01146_),
    .Q(\timer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _30532_ (.CLK(clknet_leaf_110_clk),
    .D(_01147_),
    .Q(\timer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _30533_ (.CLK(clknet_leaf_114_clk),
    .D(_01148_),
    .Q(\timer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _30534_ (.CLK(clknet_leaf_114_clk),
    .D(_01149_),
    .Q(\timer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _30535_ (.CLK(clknet_leaf_114_clk),
    .D(_01150_),
    .Q(\timer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _30536_ (.CLK(clknet_leaf_112_clk),
    .D(_01151_),
    .Q(\timer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _30537_ (.CLK(clknet_leaf_114_clk),
    .D(_01152_),
    .Q(\timer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _30538_ (.CLK(clknet_leaf_113_clk),
    .D(_01153_),
    .Q(\timer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _30539_ (.CLK(clknet_leaf_114_clk),
    .D(_01154_),
    .Q(\timer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _30540_ (.CLK(clknet_leaf_113_clk),
    .D(_01155_),
    .Q(\timer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _30541_ (.CLK(clknet_leaf_112_clk),
    .D(_01156_),
    .Q(\timer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _30542_ (.CLK(clknet_leaf_113_clk),
    .D(_01157_),
    .Q(\timer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _30543_ (.CLK(clknet_leaf_113_clk),
    .D(_01158_),
    .Q(\timer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _30544_ (.CLK(clknet_leaf_76_clk),
    .D(_01159_),
    .Q(\timer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _30545_ (.CLK(clknet_leaf_75_clk),
    .D(_01160_),
    .Q(\timer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _30546_ (.CLK(clknet_leaf_75_clk),
    .D(_01161_),
    .Q(\timer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _30547_ (.CLK(clknet_leaf_113_clk),
    .D(_01162_),
    .Q(\timer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _30548_ (.CLK(clknet_leaf_76_clk),
    .D(_01163_),
    .Q(\timer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _30549_ (.CLK(clknet_leaf_95_clk),
    .D(_01164_),
    .Q(\irq_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30550_ (.CLK(clknet_leaf_90_clk),
    .D(_01165_),
    .Q(\irq_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30551_ (.CLK(clknet_leaf_90_clk),
    .D(_01166_),
    .Q(latched_store));
 sky130_fd_sc_hd__dfxtp_1 _30552_ (.CLK(clknet_leaf_89_clk),
    .D(_01167_),
    .Q(latched_stalu));
 sky130_fd_sc_hd__dfxtp_1 _30553_ (.CLK(clknet_leaf_90_clk),
    .D(_01168_),
    .Q(latched_branch));
 sky130_fd_sc_hd__dfxtp_1 _30554_ (.CLK(clknet_leaf_90_clk),
    .D(_01169_),
    .Q(decoder_pseudo_trigger));
 sky130_fd_sc_hd__dfxtp_1 _30555_ (.CLK(clknet_leaf_85_clk),
    .D(_01170_),
    .Q(latched_is_lh));
 sky130_fd_sc_hd__dfxtp_1 _30556_ (.CLK(clknet_leaf_85_clk),
    .D(_01171_),
    .Q(latched_is_lb));
 sky130_fd_sc_hd__dfxtp_1 _30557_ (.CLK(clknet_leaf_52_clk),
    .D(_01172_),
    .Q(\pcpi_timeout_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30558_ (.CLK(clknet_leaf_51_clk),
    .D(_01173_),
    .Q(\pcpi_timeout_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30559_ (.CLK(clknet_leaf_52_clk),
    .D(_01174_),
    .Q(\pcpi_timeout_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30560_ (.CLK(clknet_leaf_52_clk),
    .D(_01175_),
    .Q(\pcpi_timeout_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30561_ (.CLK(clknet_leaf_63_clk),
    .D(_01176_),
    .Q(pcpi_timeout));
 sky130_fd_sc_hd__dfxtp_1 _30562_ (.CLK(clknet_leaf_34_clk),
    .D(\alu_out[0] ),
    .Q(\alu_out_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30563_ (.CLK(clknet_leaf_34_clk),
    .D(\alu_out[1] ),
    .Q(\alu_out_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30564_ (.CLK(clknet_leaf_47_clk),
    .D(\alu_out[2] ),
    .Q(\alu_out_q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30565_ (.CLK(clknet_leaf_34_clk),
    .D(\alu_out[3] ),
    .Q(\alu_out_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30566_ (.CLK(clknet_leaf_34_clk),
    .D(\alu_out[4] ),
    .Q(\alu_out_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _30567_ (.CLK(clknet_leaf_34_clk),
    .D(\alu_out[5] ),
    .Q(\alu_out_q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _30568_ (.CLK(clknet_leaf_35_clk),
    .D(\alu_out[6] ),
    .Q(\alu_out_q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _30569_ (.CLK(clknet_leaf_35_clk),
    .D(\alu_out[7] ),
    .Q(\alu_out_q[7] ));
 sky130_fd_sc_hd__dfxtp_1 _30570_ (.CLK(clknet_leaf_35_clk),
    .D(\alu_out[8] ),
    .Q(\alu_out_q[8] ));
 sky130_fd_sc_hd__dfxtp_1 _30571_ (.CLK(clknet_leaf_35_clk),
    .D(\alu_out[9] ),
    .Q(\alu_out_q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _30572_ (.CLK(clknet_leaf_36_clk),
    .D(\alu_out[10] ),
    .Q(\alu_out_q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _30573_ (.CLK(clknet_leaf_36_clk),
    .D(\alu_out[11] ),
    .Q(\alu_out_q[11] ));
 sky130_fd_sc_hd__dfxtp_1 _30574_ (.CLK(clknet_leaf_36_clk),
    .D(\alu_out[12] ),
    .Q(\alu_out_q[12] ));
 sky130_fd_sc_hd__dfxtp_1 _30575_ (.CLK(clknet_leaf_12_clk),
    .D(\alu_out[13] ),
    .Q(\alu_out_q[13] ));
 sky130_fd_sc_hd__dfxtp_1 _30576_ (.CLK(clknet_leaf_20_clk),
    .D(\alu_out[14] ),
    .Q(\alu_out_q[14] ));
 sky130_fd_sc_hd__dfxtp_1 _30577_ (.CLK(clknet_leaf_19_clk),
    .D(\alu_out[15] ),
    .Q(\alu_out_q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _30578_ (.CLK(clknet_leaf_13_clk),
    .D(\alu_out[16] ),
    .Q(\alu_out_q[16] ));
 sky130_fd_sc_hd__dfxtp_1 _30579_ (.CLK(clknet_leaf_15_clk),
    .D(\alu_out[17] ),
    .Q(\alu_out_q[17] ));
 sky130_fd_sc_hd__dfxtp_1 _30580_ (.CLK(clknet_leaf_18_clk),
    .D(\alu_out[18] ),
    .Q(\alu_out_q[18] ));
 sky130_fd_sc_hd__dfxtp_1 _30581_ (.CLK(clknet_leaf_212_clk),
    .D(\alu_out[19] ),
    .Q(\alu_out_q[19] ));
 sky130_fd_sc_hd__dfxtp_1 _30582_ (.CLK(clknet_leaf_17_clk),
    .D(\alu_out[20] ),
    .Q(\alu_out_q[20] ));
 sky130_fd_sc_hd__dfxtp_1 _30583_ (.CLK(clknet_leaf_18_clk),
    .D(\alu_out[21] ),
    .Q(\alu_out_q[21] ));
 sky130_fd_sc_hd__dfxtp_1 _30584_ (.CLK(clknet_leaf_17_clk),
    .D(\alu_out[22] ),
    .Q(\alu_out_q[22] ));
 sky130_fd_sc_hd__dfxtp_1 _30585_ (.CLK(clknet_leaf_211_clk),
    .D(\alu_out[23] ),
    .Q(\alu_out_q[23] ));
 sky130_fd_sc_hd__dfxtp_1 _30586_ (.CLK(clknet_leaf_15_clk),
    .D(\alu_out[24] ),
    .Q(\alu_out_q[24] ));
 sky130_fd_sc_hd__dfxtp_1 _30587_ (.CLK(clknet_leaf_15_clk),
    .D(\alu_out[25] ),
    .Q(\alu_out_q[25] ));
 sky130_fd_sc_hd__dfxtp_1 _30588_ (.CLK(clknet_leaf_17_clk),
    .D(\alu_out[26] ),
    .Q(\alu_out_q[26] ));
 sky130_fd_sc_hd__dfxtp_1 _30589_ (.CLK(clknet_leaf_209_clk),
    .D(\alu_out[27] ),
    .Q(\alu_out_q[27] ));
 sky130_fd_sc_hd__dfxtp_1 _30590_ (.CLK(clknet_leaf_13_clk),
    .D(net423),
    .Q(\alu_out_q[28] ));
 sky130_fd_sc_hd__dfxtp_1 _30591_ (.CLK(clknet_leaf_209_clk),
    .D(\alu_out[29] ),
    .Q(\alu_out_q[29] ));
 sky130_fd_sc_hd__dfxtp_1 _30592_ (.CLK(clknet_leaf_21_clk),
    .D(\alu_out[30] ),
    .Q(\alu_out_q[30] ));
 sky130_fd_sc_hd__dfxtp_1 _30593_ (.CLK(clknet_leaf_12_clk),
    .D(\alu_out[31] ),
    .Q(\alu_out_q[31] ));
 sky130_fd_sc_hd__dfxtp_1 _30594_ (.CLK(clknet_leaf_95_clk),
    .D(_01177_),
    .Q(do_waitirq));
 sky130_fd_sc_hd__dfxtp_1 _30595_ (.CLK(clknet_leaf_66_clk),
    .D(_01178_),
    .Q(net235));
 sky130_fd_sc_hd__dfxtp_1 _30596_ (.CLK(clknet_leaf_66_clk),
    .D(_01179_),
    .Q(net246));
 sky130_fd_sc_hd__dfxtp_1 _30597_ (.CLK(clknet_leaf_66_clk),
    .D(_01180_),
    .Q(net257));
 sky130_fd_sc_hd__dfxtp_1 _30598_ (.CLK(clknet_leaf_65_clk),
    .D(_01181_),
    .Q(net260));
 sky130_fd_sc_hd__dfxtp_1 _30599_ (.CLK(clknet_leaf_63_clk),
    .D(_01182_),
    .Q(net261));
 sky130_fd_sc_hd__dfxtp_1 _30600_ (.CLK(clknet_leaf_63_clk),
    .D(_01183_),
    .Q(net262));
 sky130_fd_sc_hd__dfxtp_1 _30601_ (.CLK(clknet_leaf_65_clk),
    .D(_01184_),
    .Q(net263));
 sky130_fd_sc_hd__dfxtp_1 _30602_ (.CLK(clknet_leaf_67_clk),
    .D(_01185_),
    .Q(net264));
 sky130_fd_sc_hd__dfxtp_1 _30603_ (.CLK(clknet_leaf_71_clk),
    .D(_01186_),
    .Q(net265));
 sky130_fd_sc_hd__dfxtp_1 _30604_ (.CLK(clknet_leaf_71_clk),
    .D(_01187_),
    .Q(net266));
 sky130_fd_sc_hd__dfxtp_1 _30605_ (.CLK(clknet_leaf_71_clk),
    .D(_01188_),
    .Q(net236));
 sky130_fd_sc_hd__dfxtp_1 _30606_ (.CLK(clknet_leaf_74_clk),
    .D(_01189_),
    .Q(net237));
 sky130_fd_sc_hd__dfxtp_2 _30607_ (.CLK(clknet_leaf_12_clk),
    .D(_01190_),
    .Q(net238));
 sky130_fd_sc_hd__dfxtp_2 _30608_ (.CLK(clknet_leaf_20_clk),
    .D(_01191_),
    .Q(net239));
 sky130_fd_sc_hd__dfxtp_2 _30609_ (.CLK(clknet_leaf_49_clk),
    .D(_01192_),
    .Q(net240));
 sky130_fd_sc_hd__dfxtp_1 _30610_ (.CLK(clknet_leaf_73_clk),
    .D(_01193_),
    .Q(net241));
 sky130_fd_sc_hd__dfxtp_1 _30611_ (.CLK(clknet_leaf_74_clk),
    .D(_01194_),
    .Q(net242));
 sky130_fd_sc_hd__dfxtp_1 _30612_ (.CLK(clknet_leaf_74_clk),
    .D(_01195_),
    .Q(net243));
 sky130_fd_sc_hd__dfxtp_1 _30613_ (.CLK(clknet_leaf_74_clk),
    .D(_01196_),
    .Q(net244));
 sky130_fd_sc_hd__dfxtp_1 _30614_ (.CLK(clknet_leaf_74_clk),
    .D(_01197_),
    .Q(net245));
 sky130_fd_sc_hd__dfxtp_1 _30615_ (.CLK(clknet_leaf_71_clk),
    .D(_01198_),
    .Q(net247));
 sky130_fd_sc_hd__dfxtp_1 _30616_ (.CLK(clknet_leaf_70_clk),
    .D(_01199_),
    .Q(net248));
 sky130_fd_sc_hd__dfxtp_1 _30617_ (.CLK(clknet_leaf_71_clk),
    .D(_01200_),
    .Q(net249));
 sky130_fd_sc_hd__dfxtp_2 _30618_ (.CLK(clknet_leaf_32_clk),
    .D(_01201_),
    .Q(net250));
 sky130_fd_sc_hd__dfxtp_1 _30619_ (.CLK(clknet_leaf_33_clk),
    .D(_01202_),
    .Q(net251));
 sky130_fd_sc_hd__dfxtp_2 _30620_ (.CLK(clknet_leaf_64_clk),
    .D(_01203_),
    .Q(net252));
 sky130_fd_sc_hd__dfxtp_2 _30621_ (.CLK(clknet_leaf_63_clk),
    .D(_01204_),
    .Q(net253));
 sky130_fd_sc_hd__dfxtp_1 _30622_ (.CLK(clknet_leaf_64_clk),
    .D(_01205_),
    .Q(net254));
 sky130_fd_sc_hd__dfxtp_2 _30623_ (.CLK(clknet_leaf_86_clk),
    .D(_01206_),
    .Q(net255));
 sky130_fd_sc_hd__dfxtp_1 _30624_ (.CLK(clknet_leaf_32_clk),
    .D(_01207_),
    .Q(net256));
 sky130_fd_sc_hd__dfxtp_2 _30625_ (.CLK(clknet_leaf_32_clk),
    .D(_01208_),
    .Q(net258));
 sky130_fd_sc_hd__dfxtp_1 _30626_ (.CLK(clknet_leaf_49_clk),
    .D(_01209_),
    .Q(net259));
 sky130_fd_sc_hd__dfxtp_1 _30627_ (.CLK(clknet_leaf_86_clk),
    .D(_01210_),
    .Q(instr_lui));
 sky130_fd_sc_hd__dfxtp_1 _30628_ (.CLK(clknet_leaf_86_clk),
    .D(_01211_),
    .Q(instr_auipc));
 sky130_fd_sc_hd__dfxtp_1 _30629_ (.CLK(clknet_leaf_30_clk),
    .D(_01212_),
    .Q(instr_jal));
 sky130_fd_sc_hd__dfxtp_1 _30630_ (.CLK(clknet_leaf_52_clk),
    .D(_01213_),
    .Q(instr_beq));
 sky130_fd_sc_hd__dfxtp_1 _30631_ (.CLK(clknet_leaf_51_clk),
    .D(_01214_),
    .Q(instr_bne));
 sky130_fd_sc_hd__dfxtp_1 _30632_ (.CLK(clknet_leaf_52_clk),
    .D(_01215_),
    .Q(instr_blt));
 sky130_fd_sc_hd__dfxtp_1 _30633_ (.CLK(clknet_leaf_48_clk),
    .D(_01216_),
    .Q(instr_bge));
 sky130_fd_sc_hd__dfxtp_1 _30634_ (.CLK(clknet_leaf_45_clk),
    .D(_01217_),
    .Q(instr_bltu));
 sky130_fd_sc_hd__dfxtp_1 _30635_ (.CLK(clknet_leaf_48_clk),
    .D(_01218_),
    .Q(instr_bgeu));
 sky130_fd_sc_hd__dfxtp_2 _30636_ (.CLK(clknet_leaf_87_clk),
    .D(_01219_),
    .Q(instr_jalr));
 sky130_fd_sc_hd__dfxtp_1 _30637_ (.CLK(clknet_leaf_50_clk),
    .D(_01220_),
    .Q(instr_lb));
 sky130_fd_sc_hd__dfxtp_1 _30638_ (.CLK(clknet_leaf_50_clk),
    .D(_01221_),
    .Q(instr_lh));
 sky130_fd_sc_hd__dfxtp_1 _30639_ (.CLK(clknet_leaf_50_clk),
    .D(_01222_),
    .Q(instr_lw));
 sky130_fd_sc_hd__dfxtp_1 _30640_ (.CLK(clknet_leaf_50_clk),
    .D(_01223_),
    .Q(instr_lbu));
 sky130_fd_sc_hd__dfxtp_1 _30641_ (.CLK(clknet_leaf_50_clk),
    .D(_01224_),
    .Q(instr_lhu));
 sky130_fd_sc_hd__dfxtp_1 _30642_ (.CLK(clknet_leaf_50_clk),
    .D(_01225_),
    .Q(instr_sb));
 sky130_fd_sc_hd__dfxtp_1 _30643_ (.CLK(clknet_leaf_49_clk),
    .D(_01226_),
    .Q(instr_sh));
 sky130_fd_sc_hd__dfxtp_1 _30644_ (.CLK(clknet_leaf_50_clk),
    .D(_01227_),
    .Q(instr_addi));
 sky130_fd_sc_hd__dfxtp_1 _30645_ (.CLK(clknet_leaf_53_clk),
    .D(_01228_),
    .Q(instr_slti));
 sky130_fd_sc_hd__dfxtp_1 _30646_ (.CLK(clknet_leaf_53_clk),
    .D(_01229_),
    .Q(instr_sltiu));
 sky130_fd_sc_hd__dfxtp_1 _30647_ (.CLK(clknet_leaf_53_clk),
    .D(_01230_),
    .Q(instr_xori));
 sky130_fd_sc_hd__dfxtp_1 _30648_ (.CLK(clknet_leaf_44_clk),
    .D(_01231_),
    .Q(instr_ori));
 sky130_fd_sc_hd__dfxtp_1 _30649_ (.CLK(clknet_leaf_45_clk),
    .D(_01232_),
    .Q(instr_andi));
 sky130_fd_sc_hd__dfxtp_1 _30650_ (.CLK(clknet_leaf_63_clk),
    .D(_01233_),
    .Q(instr_sw));
 sky130_fd_sc_hd__dfxtp_1 _30651_ (.CLK(clknet_leaf_49_clk),
    .D(_01234_),
    .Q(instr_slli));
 sky130_fd_sc_hd__dfxtp_1 _30652_ (.CLK(clknet_leaf_51_clk),
    .D(_01235_),
    .Q(instr_srli));
 sky130_fd_sc_hd__dfxtp_1 _30653_ (.CLK(clknet_leaf_50_clk),
    .D(_01236_),
    .Q(instr_add));
 sky130_fd_sc_hd__dfxtp_2 _30654_ (.CLK(clknet_leaf_48_clk),
    .D(_01237_),
    .Q(instr_sub));
 sky130_fd_sc_hd__dfxtp_1 _30655_ (.CLK(clknet_leaf_51_clk),
    .D(_01238_),
    .Q(instr_sll));
 sky130_fd_sc_hd__dfxtp_1 _30656_ (.CLK(clknet_leaf_52_clk),
    .D(_01239_),
    .Q(instr_slt));
 sky130_fd_sc_hd__dfxtp_1 _30657_ (.CLK(clknet_leaf_44_clk),
    .D(_01240_),
    .Q(instr_sltu));
 sky130_fd_sc_hd__dfxtp_1 _30658_ (.CLK(clknet_leaf_51_clk),
    .D(_01241_),
    .Q(instr_xor));
 sky130_fd_sc_hd__dfxtp_1 _30659_ (.CLK(clknet_leaf_50_clk),
    .D(_01242_),
    .Q(instr_srl));
 sky130_fd_sc_hd__dfxtp_2 _30660_ (.CLK(clknet_leaf_48_clk),
    .D(_01243_),
    .Q(instr_sra));
 sky130_fd_sc_hd__dfxtp_1 _30661_ (.CLK(clknet_leaf_45_clk),
    .D(_01244_),
    .Q(instr_or));
 sky130_fd_sc_hd__dfxtp_1 _30662_ (.CLK(clknet_leaf_48_clk),
    .D(_01245_),
    .Q(instr_and));
 sky130_fd_sc_hd__dfxtp_2 _30663_ (.CLK(clknet_leaf_48_clk),
    .D(_01246_),
    .Q(instr_srai));
 sky130_fd_sc_hd__dfxtp_1 _30664_ (.CLK(clknet_leaf_66_clk),
    .D(_01247_),
    .Q(instr_rdcycle));
 sky130_fd_sc_hd__dfxtp_1 _30665_ (.CLK(clknet_leaf_66_clk),
    .D(_01248_),
    .Q(instr_rdcycleh));
 sky130_fd_sc_hd__dfxtp_1 _30666_ (.CLK(clknet_leaf_68_clk),
    .D(_01249_),
    .Q(instr_rdinstr));
 sky130_fd_sc_hd__dfxtp_1 _30667_ (.CLK(clknet_leaf_68_clk),
    .D(_01250_),
    .Q(instr_rdinstrh));
 sky130_fd_sc_hd__dfxtp_1 _30668_ (.CLK(clknet_leaf_65_clk),
    .D(_01251_),
    .Q(instr_ecall_ebreak));
 sky130_fd_sc_hd__dfxtp_1 _30669_ (.CLK(clknet_leaf_67_clk),
    .D(_01252_),
    .Q(instr_getq));
 sky130_fd_sc_hd__dfxtp_2 _30670_ (.CLK(clknet_leaf_67_clk),
    .D(_01253_),
    .Q(instr_setq));
 sky130_fd_sc_hd__dfxtp_1 _30671_ (.CLK(clknet_leaf_89_clk),
    .D(_01254_),
    .Q(instr_retirq));
 sky130_fd_sc_hd__dfxtp_1 _30672_ (.CLK(clknet_leaf_72_clk),
    .D(_01255_),
    .Q(instr_maskirq));
 sky130_fd_sc_hd__dfxtp_1 _30673_ (.CLK(clknet_leaf_95_clk),
    .D(_01256_),
    .Q(instr_waitirq));
 sky130_fd_sc_hd__dfxtp_1 _30674_ (.CLK(clknet_leaf_67_clk),
    .D(_01257_),
    .Q(instr_timer));
 sky130_fd_sc_hd__dfxtp_1 _30675_ (.CLK(clknet_leaf_97_clk),
    .D(_01258_),
    .Q(\decoded_rs1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30676_ (.CLK(clknet_leaf_97_clk),
    .D(_01259_),
    .Q(\decoded_rs1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30677_ (.CLK(clknet_leaf_96_clk),
    .D(_01260_),
    .Q(\decoded_rs1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30678_ (.CLK(clknet_leaf_96_clk),
    .D(_01261_),
    .Q(\decoded_rs1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30679_ (.CLK(clknet_leaf_104_clk),
    .D(_01262_),
    .Q(\decoded_rd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30680_ (.CLK(clknet_leaf_105_clk),
    .D(_01263_),
    .Q(\decoded_rd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30681_ (.CLK(clknet_leaf_104_clk),
    .D(_01264_),
    .Q(\decoded_rd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30682_ (.CLK(clknet_leaf_109_clk),
    .D(_01265_),
    .Q(\decoded_rd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30683_ (.CLK(clknet_leaf_97_clk),
    .D(_01266_),
    .Q(\decoded_rd[4] ));
 sky130_fd_sc_hd__dfxtp_1 _30684_ (.CLK(clknet_leaf_29_clk),
    .D(_01267_),
    .Q(\decoded_imm_uj[11] ));
 sky130_fd_sc_hd__dfxtp_1 _30685_ (.CLK(clknet_leaf_95_clk),
    .D(_01268_),
    .Q(\decoded_imm_uj[1] ));
 sky130_fd_sc_hd__dfxtp_2 _30686_ (.CLK(clknet_leaf_33_clk),
    .D(_01269_),
    .Q(\decoded_imm_uj[2] ));
 sky130_fd_sc_hd__dfxtp_2 _30687_ (.CLK(clknet_leaf_31_clk),
    .D(_01270_),
    .Q(\decoded_imm_uj[3] ));
 sky130_fd_sc_hd__dfxtp_2 _30688_ (.CLK(clknet_leaf_30_clk),
    .D(_01271_),
    .Q(\decoded_imm[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30689_ (.CLK(clknet_leaf_24_clk),
    .D(_00037_),
    .Q(is_lui_auipc_jal));
 sky130_fd_sc_hd__dfxtp_1 _30690_ (.CLK(clknet_leaf_85_clk),
    .D(_01272_),
    .Q(is_lb_lh_lw_lbu_lhu));
 sky130_fd_sc_hd__dfxtp_1 _30691_ (.CLK(clknet_leaf_32_clk),
    .D(_01273_),
    .Q(is_slli_srli_srai));
 sky130_fd_sc_hd__dfxtp_1 _30692_ (.CLK(clknet_leaf_87_clk),
    .D(_01274_),
    .Q(is_jalr_addi_slti_sltiu_xori_ori_andi));
 sky130_fd_sc_hd__dfxtp_1 _30693_ (.CLK(clknet_leaf_85_clk),
    .D(_01275_),
    .Q(is_sb_sh_sw));
 sky130_fd_sc_hd__dfxtp_1 _30694_ (.CLK(clknet_leaf_45_clk),
    .D(_00038_),
    .Q(is_slti_blt_slt));
 sky130_fd_sc_hd__dfxtp_1 _30695_ (.CLK(clknet_leaf_45_clk),
    .D(_00039_),
    .Q(is_sltiu_bltu_sltu));
 sky130_fd_sc_hd__dfxtp_1 _30696_ (.CLK(clknet_leaf_85_clk),
    .D(_01276_),
    .Q(is_beq_bne_blt_bge_bltu_bgeu));
 sky130_fd_sc_hd__dfxtp_1 _30697_ (.CLK(clknet_leaf_86_clk),
    .D(_01277_),
    .Q(is_alu_reg_imm));
 sky130_fd_sc_hd__dfxtp_1 _30698_ (.CLK(clknet_leaf_86_clk),
    .D(_01278_),
    .Q(is_alu_reg_reg));
 sky130_fd_sc_hd__dfxtp_1 _30699_ (.CLK(clknet_leaf_47_clk),
    .D(_01279_),
    .Q(is_compare));
 sky130_fd_sc_hd__dfxtp_2 _30700_ (.CLK(clknet_leaf_84_clk),
    .D(_01280_),
    .Q(net129));
 sky130_fd_sc_hd__dfxtp_1 _30701_ (.CLK(clknet_leaf_83_clk),
    .D(_01281_),
    .Q(\mem_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30702_ (.CLK(clknet_leaf_67_clk),
    .D(_01282_),
    .Q(\mem_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30703_ (.CLK(clknet_leaf_44_clk),
    .D(_01283_),
    .Q(net199));
 sky130_fd_sc_hd__dfxtp_1 _30704_ (.CLK(clknet_leaf_44_clk),
    .D(_01284_),
    .Q(net210));
 sky130_fd_sc_hd__dfxtp_1 _30705_ (.CLK(clknet_leaf_42_clk),
    .D(_01285_),
    .Q(net221));
 sky130_fd_sc_hd__dfxtp_1 _30706_ (.CLK(clknet_leaf_40_clk),
    .D(_01286_),
    .Q(net224));
 sky130_fd_sc_hd__dfxtp_1 _30707_ (.CLK(clknet_leaf_43_clk),
    .D(_01287_),
    .Q(net225));
 sky130_fd_sc_hd__dfxtp_1 _30708_ (.CLK(clknet_leaf_43_clk),
    .D(_01288_),
    .Q(net226));
 sky130_fd_sc_hd__dfxtp_1 _30709_ (.CLK(clknet_leaf_43_clk),
    .D(_01289_),
    .Q(net227));
 sky130_fd_sc_hd__dfxtp_1 _30710_ (.CLK(clknet_leaf_43_clk),
    .D(_01290_),
    .Q(net228));
 sky130_fd_sc_hd__dfxtp_1 _30711_ (.CLK(clknet_leaf_42_clk),
    .D(_01291_),
    .Q(net229));
 sky130_fd_sc_hd__dfxtp_1 _30712_ (.CLK(clknet_leaf_43_clk),
    .D(_01292_),
    .Q(net230));
 sky130_fd_sc_hd__dfxtp_1 _30713_ (.CLK(clknet_leaf_42_clk),
    .D(_01293_),
    .Q(net200));
 sky130_fd_sc_hd__dfxtp_1 _30714_ (.CLK(clknet_leaf_42_clk),
    .D(_01294_),
    .Q(net201));
 sky130_fd_sc_hd__dfxtp_2 _30715_ (.CLK(clknet_leaf_42_clk),
    .D(_01295_),
    .Q(net202));
 sky130_fd_sc_hd__dfxtp_1 _30716_ (.CLK(clknet_leaf_42_clk),
    .D(_01296_),
    .Q(net203));
 sky130_fd_sc_hd__dfxtp_1 _30717_ (.CLK(clknet_leaf_45_clk),
    .D(_01297_),
    .Q(net204));
 sky130_fd_sc_hd__dfxtp_1 _30718_ (.CLK(clknet_leaf_47_clk),
    .D(_01298_),
    .Q(net205));
 sky130_fd_sc_hd__dfxtp_1 _30719_ (.CLK(clknet_leaf_40_clk),
    .D(_01299_),
    .Q(net206));
 sky130_fd_sc_hd__dfxtp_1 _30720_ (.CLK(clknet_leaf_40_clk),
    .D(_01300_),
    .Q(net207));
 sky130_fd_sc_hd__dfxtp_1 _30721_ (.CLK(clknet_leaf_42_clk),
    .D(_01301_),
    .Q(net208));
 sky130_fd_sc_hd__dfxtp_1 _30722_ (.CLK(clknet_leaf_42_clk),
    .D(_01302_),
    .Q(net209));
 sky130_fd_sc_hd__dfxtp_1 _30723_ (.CLK(clknet_leaf_3_clk),
    .D(_01303_),
    .Q(net211));
 sky130_fd_sc_hd__dfxtp_1 _30724_ (.CLK(clknet_leaf_3_clk),
    .D(_01304_),
    .Q(net212));
 sky130_fd_sc_hd__dfxtp_1 _30725_ (.CLK(clknet_leaf_3_clk),
    .D(_01305_),
    .Q(net213));
 sky130_fd_sc_hd__dfxtp_1 _30726_ (.CLK(clknet_leaf_3_clk),
    .D(_01306_),
    .Q(net214));
 sky130_fd_sc_hd__dfxtp_1 _30727_ (.CLK(clknet_leaf_42_clk),
    .D(_01307_),
    .Q(net215));
 sky130_fd_sc_hd__dfxtp_1 _30728_ (.CLK(clknet_leaf_44_clk),
    .D(_01308_),
    .Q(net216));
 sky130_fd_sc_hd__dfxtp_1 _30729_ (.CLK(clknet_leaf_46_clk),
    .D(_01309_),
    .Q(net217));
 sky130_fd_sc_hd__dfxtp_1 _30730_ (.CLK(clknet_leaf_46_clk),
    .D(_01310_),
    .Q(net218));
 sky130_fd_sc_hd__dfxtp_1 _30731_ (.CLK(clknet_leaf_47_clk),
    .D(_01311_),
    .Q(net219));
 sky130_fd_sc_hd__dfxtp_1 _30732_ (.CLK(clknet_leaf_47_clk),
    .D(_01312_),
    .Q(net220));
 sky130_fd_sc_hd__dfxtp_1 _30733_ (.CLK(clknet_leaf_47_clk),
    .D(_01313_),
    .Q(net222));
 sky130_fd_sc_hd__dfxtp_2 _30734_ (.CLK(clknet_leaf_48_clk),
    .D(_01314_),
    .Q(net223));
 sky130_fd_sc_hd__dfxtp_1 _30735_ (.CLK(clknet_leaf_45_clk),
    .D(_01315_),
    .Q(net231));
 sky130_fd_sc_hd__dfxtp_2 _30736_ (.CLK(clknet_leaf_44_clk),
    .D(_01316_),
    .Q(net232));
 sky130_fd_sc_hd__dfxtp_1 _30737_ (.CLK(clknet_leaf_44_clk),
    .D(_01317_),
    .Q(net233));
 sky130_fd_sc_hd__dfxtp_1 _30738_ (.CLK(clknet_leaf_45_clk),
    .D(_01318_),
    .Q(net234));
 sky130_fd_sc_hd__dfxtp_1 _30739_ (.CLK(clknet_leaf_47_clk),
    .D(_00000_),
    .Q(\alu_add_sub[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30740_ (.CLK(clknet_leaf_46_clk),
    .D(_00011_),
    .Q(\alu_add_sub[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30741_ (.CLK(clknet_leaf_46_clk),
    .D(_00022_),
    .Q(\alu_add_sub[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30742_ (.CLK(clknet_leaf_41_clk),
    .D(_00025_),
    .Q(\alu_add_sub[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30743_ (.CLK(clknet_leaf_47_clk),
    .D(_00026_),
    .Q(\alu_add_sub[4] ));
 sky130_fd_sc_hd__dfxtp_1 _30744_ (.CLK(clknet_leaf_34_clk),
    .D(_00027_),
    .Q(\alu_add_sub[5] ));
 sky130_fd_sc_hd__dfxtp_1 _30745_ (.CLK(clknet_leaf_35_clk),
    .D(_00028_),
    .Q(\alu_add_sub[6] ));
 sky130_fd_sc_hd__dfxtp_1 _30746_ (.CLK(clknet_leaf_37_clk),
    .D(_00029_),
    .Q(\alu_add_sub[7] ));
 sky130_fd_sc_hd__dfxtp_1 _30747_ (.CLK(clknet_leaf_38_clk),
    .D(_00030_),
    .Q(\alu_add_sub[8] ));
 sky130_fd_sc_hd__dfxtp_1 _30748_ (.CLK(clknet_leaf_37_clk),
    .D(_00031_),
    .Q(\alu_add_sub[9] ));
 sky130_fd_sc_hd__dfxtp_1 _30749_ (.CLK(clknet_leaf_37_clk),
    .D(_00001_),
    .Q(\alu_add_sub[10] ));
 sky130_fd_sc_hd__dfxtp_1 _30750_ (.CLK(clknet_leaf_11_clk),
    .D(_00002_),
    .Q(\alu_add_sub[11] ));
 sky130_fd_sc_hd__dfxtp_1 _30751_ (.CLK(clknet_leaf_36_clk),
    .D(_00003_),
    .Q(\alu_add_sub[12] ));
 sky130_fd_sc_hd__dfxtp_1 _30752_ (.CLK(clknet_leaf_12_clk),
    .D(_00004_),
    .Q(\alu_add_sub[13] ));
 sky130_fd_sc_hd__dfxtp_1 _30753_ (.CLK(clknet_leaf_11_clk),
    .D(_00005_),
    .Q(\alu_add_sub[14] ));
 sky130_fd_sc_hd__dfxtp_1 _30754_ (.CLK(clknet_leaf_10_clk),
    .D(_00006_),
    .Q(\alu_add_sub[15] ));
 sky130_fd_sc_hd__dfxtp_1 _30755_ (.CLK(clknet_leaf_14_clk),
    .D(_00007_),
    .Q(\alu_add_sub[16] ));
 sky130_fd_sc_hd__dfxtp_1 _30756_ (.CLK(clknet_leaf_1_clk),
    .D(_00008_),
    .Q(\alu_add_sub[17] ));
 sky130_fd_sc_hd__dfxtp_1 _30757_ (.CLK(clknet_leaf_1_clk),
    .D(_00009_),
    .Q(\alu_add_sub[18] ));
 sky130_fd_sc_hd__dfxtp_1 _30758_ (.CLK(clknet_leaf_1_clk),
    .D(_00010_),
    .Q(\alu_add_sub[19] ));
 sky130_fd_sc_hd__dfxtp_1 _30759_ (.CLK(clknet_leaf_2_clk),
    .D(_00012_),
    .Q(\alu_add_sub[20] ));
 sky130_fd_sc_hd__dfxtp_1 _30760_ (.CLK(clknet_leaf_0_clk),
    .D(_00013_),
    .Q(\alu_add_sub[21] ));
 sky130_fd_sc_hd__dfxtp_1 _30761_ (.CLK(clknet_leaf_0_clk),
    .D(_00014_),
    .Q(\alu_add_sub[22] ));
 sky130_fd_sc_hd__dfxtp_1 _30762_ (.CLK(clknet_leaf_225_clk),
    .D(_00015_),
    .Q(\alu_add_sub[23] ));
 sky130_fd_sc_hd__dfxtp_1 _30763_ (.CLK(clknet_leaf_225_clk),
    .D(_00016_),
    .Q(\alu_add_sub[24] ));
 sky130_fd_sc_hd__dfxtp_1 _30764_ (.CLK(clknet_leaf_14_clk),
    .D(_00017_),
    .Q(\alu_add_sub[25] ));
 sky130_fd_sc_hd__dfxtp_1 _30765_ (.CLK(clknet_leaf_15_clk),
    .D(_00018_),
    .Q(\alu_add_sub[26] ));
 sky130_fd_sc_hd__dfxtp_1 _30766_ (.CLK(clknet_leaf_14_clk),
    .D(_00019_),
    .Q(\alu_add_sub[27] ));
 sky130_fd_sc_hd__dfxtp_1 _30767_ (.CLK(clknet_leaf_14_clk),
    .D(_00020_),
    .Q(\alu_add_sub[28] ));
 sky130_fd_sc_hd__dfxtp_1 _30768_ (.CLK(clknet_leaf_14_clk),
    .D(_00021_),
    .Q(\alu_add_sub[29] ));
 sky130_fd_sc_hd__dfxtp_1 _30769_ (.CLK(clknet_leaf_13_clk),
    .D(_00023_),
    .Q(\alu_add_sub[30] ));
 sky130_fd_sc_hd__dfxtp_1 _30770_ (.CLK(clknet_leaf_12_clk),
    .D(_00024_),
    .Q(\alu_add_sub[31] ));
 sky130_fd_sc_hd__dfxtp_1 _30771_ (.CLK(clknet_leaf_10_clk),
    .D(_14604_),
    .Q(\alu_shl[16] ));
 sky130_fd_sc_hd__dfxtp_1 _30772_ (.CLK(clknet_leaf_10_clk),
    .D(_14605_),
    .Q(\alu_shl[17] ));
 sky130_fd_sc_hd__dfxtp_1 _30773_ (.CLK(clknet_leaf_5_clk),
    .D(_14606_),
    .Q(\alu_shl[18] ));
 sky130_fd_sc_hd__dfxtp_1 _30774_ (.CLK(clknet_leaf_2_clk),
    .D(_14607_),
    .Q(\alu_shl[19] ));
 sky130_fd_sc_hd__dfxtp_1 _30775_ (.CLK(clknet_leaf_3_clk),
    .D(_14608_),
    .Q(\alu_shl[20] ));
 sky130_fd_sc_hd__dfxtp_1 _30776_ (.CLK(clknet_leaf_2_clk),
    .D(_14609_),
    .Q(\alu_shl[21] ));
 sky130_fd_sc_hd__dfxtp_1 _30777_ (.CLK(clknet_leaf_3_clk),
    .D(_14610_),
    .Q(\alu_shl[22] ));
 sky130_fd_sc_hd__dfxtp_1 _30778_ (.CLK(clknet_leaf_2_clk),
    .D(_14611_),
    .Q(\alu_shl[23] ));
 sky130_fd_sc_hd__dfxtp_1 _30779_ (.CLK(clknet_leaf_2_clk),
    .D(_14612_),
    .Q(\alu_shl[24] ));
 sky130_fd_sc_hd__dfxtp_1 _30780_ (.CLK(clknet_leaf_1_clk),
    .D(_14613_),
    .Q(\alu_shl[25] ));
 sky130_fd_sc_hd__dfxtp_1 _30781_ (.CLK(clknet_leaf_5_clk),
    .D(_14614_),
    .Q(\alu_shl[26] ));
 sky130_fd_sc_hd__dfxtp_1 _30782_ (.CLK(clknet_leaf_10_clk),
    .D(_14615_),
    .Q(\alu_shl[27] ));
 sky130_fd_sc_hd__dfxtp_1 _30783_ (.CLK(clknet_5_2__leaf_clk),
    .D(_14616_),
    .Q(\alu_shl[28] ));
 sky130_fd_sc_hd__dfxtp_1 _30784_ (.CLK(clknet_leaf_10_clk),
    .D(_14617_),
    .Q(\alu_shl[29] ));
 sky130_fd_sc_hd__dfxtp_1 _30785_ (.CLK(clknet_leaf_9_clk),
    .D(_14618_),
    .Q(\alu_shl[30] ));
 sky130_fd_sc_hd__dfxtp_1 _30786_ (.CLK(clknet_leaf_10_clk),
    .D(_14619_),
    .Q(\alu_shl[31] ));
 sky130_fd_sc_hd__dfxtp_1 _30787_ (.CLK(clknet_leaf_40_clk),
    .D(_14620_),
    .Q(\alu_shr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30788_ (.CLK(clknet_leaf_40_clk),
    .D(_14631_),
    .Q(\alu_shr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30789_ (.CLK(clknet_leaf_40_clk),
    .D(_14642_),
    .Q(\alu_shr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30790_ (.CLK(clknet_leaf_40_clk),
    .D(_14645_),
    .Q(\alu_shr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30791_ (.CLK(clknet_leaf_40_clk),
    .D(_14646_),
    .Q(\alu_shr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _30792_ (.CLK(clknet_leaf_40_clk),
    .D(_14647_),
    .Q(\alu_shr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _30793_ (.CLK(clknet_leaf_40_clk),
    .D(_14648_),
    .Q(\alu_shr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _30794_ (.CLK(clknet_leaf_39_clk),
    .D(_14649_),
    .Q(\alu_shr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _30795_ (.CLK(clknet_leaf_39_clk),
    .D(_14650_),
    .Q(\alu_shr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _30796_ (.CLK(clknet_leaf_38_clk),
    .D(_14651_),
    .Q(\alu_shr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _30797_ (.CLK(clknet_leaf_38_clk),
    .D(_14621_),
    .Q(\alu_shr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _30798_ (.CLK(clknet_leaf_39_clk),
    .D(_14622_),
    .Q(\alu_shr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _30799_ (.CLK(clknet_leaf_39_clk),
    .D(_14623_),
    .Q(\alu_shr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _30800_ (.CLK(clknet_leaf_8_clk),
    .D(_14624_),
    .Q(\alu_shr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _30801_ (.CLK(clknet_leaf_9_clk),
    .D(_14625_),
    .Q(\alu_shr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _30802_ (.CLK(clknet_leaf_8_clk),
    .D(_14626_),
    .Q(\alu_shr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _30803_ (.CLK(clknet_leaf_5_clk),
    .D(_14627_),
    .Q(\alu_shr[16] ));
 sky130_fd_sc_hd__dfxtp_1 _30804_ (.CLK(clknet_leaf_5_clk),
    .D(_14628_),
    .Q(\alu_shr[17] ));
 sky130_fd_sc_hd__dfxtp_1 _30805_ (.CLK(clknet_leaf_5_clk),
    .D(_14629_),
    .Q(\alu_shr[18] ));
 sky130_fd_sc_hd__dfxtp_1 _30806_ (.CLK(clknet_leaf_5_clk),
    .D(_14630_),
    .Q(\alu_shr[19] ));
 sky130_fd_sc_hd__dfxtp_1 _30807_ (.CLK(clknet_leaf_5_clk),
    .D(_14632_),
    .Q(\alu_shr[20] ));
 sky130_fd_sc_hd__dfxtp_1 _30808_ (.CLK(clknet_leaf_4_clk),
    .D(_14633_),
    .Q(\alu_shr[21] ));
 sky130_fd_sc_hd__dfxtp_1 _30809_ (.CLK(clknet_leaf_4_clk),
    .D(_14634_),
    .Q(\alu_shr[22] ));
 sky130_fd_sc_hd__dfxtp_1 _30810_ (.CLK(clknet_leaf_5_clk),
    .D(_14635_),
    .Q(\alu_shr[23] ));
 sky130_fd_sc_hd__dfxtp_1 _30811_ (.CLK(clknet_leaf_5_clk),
    .D(_14636_),
    .Q(\alu_shr[24] ));
 sky130_fd_sc_hd__dfxtp_1 _30812_ (.CLK(clknet_leaf_5_clk),
    .D(_14637_),
    .Q(\alu_shr[25] ));
 sky130_fd_sc_hd__dfxtp_1 _30813_ (.CLK(clknet_leaf_5_clk),
    .D(_14638_),
    .Q(\alu_shr[26] ));
 sky130_fd_sc_hd__dfxtp_1 _30814_ (.CLK(clknet_leaf_5_clk),
    .D(_14639_),
    .Q(\alu_shr[27] ));
 sky130_fd_sc_hd__dfxtp_1 _30815_ (.CLK(clknet_5_2__leaf_clk),
    .D(_14640_),
    .Q(\alu_shr[28] ));
 sky130_fd_sc_hd__dfxtp_1 _30816_ (.CLK(clknet_leaf_8_clk),
    .D(_14641_),
    .Q(\alu_shr[29] ));
 sky130_fd_sc_hd__dfxtp_1 _30817_ (.CLK(clknet_leaf_8_clk),
    .D(_14643_),
    .Q(\alu_shr[30] ));
 sky130_fd_sc_hd__dfxtp_1 _30818_ (.CLK(clknet_leaf_9_clk),
    .D(_14644_),
    .Q(\alu_shr[31] ));
 sky130_fd_sc_hd__dfxtp_1 _30819_ (.CLK(clknet_leaf_47_clk),
    .D(_00032_),
    .Q(alu_eq));
 sky130_fd_sc_hd__dfxtp_1 _30820_ (.CLK(clknet_leaf_47_clk),
    .D(_00034_),
    .Q(alu_ltu));
 sky130_fd_sc_hd__dfxtp_1 _30821_ (.CLK(clknet_leaf_48_clk),
    .D(_00033_),
    .Q(alu_lts));
 sky130_fd_sc_hd__dfxtp_1 _30822_ (.CLK(clknet_leaf_38_clk),
    .D(_01319_),
    .Q(\alu_shl[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30823_ (.CLK(clknet_leaf_41_clk),
    .D(_01320_),
    .Q(\alu_shl[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30824_ (.CLK(clknet_leaf_40_clk),
    .D(_01321_),
    .Q(\alu_shl[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30825_ (.CLK(clknet_leaf_41_clk),
    .D(_01322_),
    .Q(\alu_shl[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30826_ (.CLK(clknet_leaf_40_clk),
    .D(_01323_),
    .Q(\alu_shl[4] ));
 sky130_fd_sc_hd__dfxtp_1 _30827_ (.CLK(clknet_leaf_38_clk),
    .D(_01324_),
    .Q(\alu_shl[5] ));
 sky130_fd_sc_hd__dfxtp_1 _30828_ (.CLK(clknet_leaf_40_clk),
    .D(_01325_),
    .Q(\alu_shl[6] ));
 sky130_fd_sc_hd__dfxtp_1 _30829_ (.CLK(clknet_leaf_38_clk),
    .D(_01326_),
    .Q(\alu_shl[7] ));
 sky130_fd_sc_hd__dfxtp_1 _30830_ (.CLK(clknet_leaf_38_clk),
    .D(_01327_),
    .Q(\alu_shl[8] ));
 sky130_fd_sc_hd__dfxtp_1 _30831_ (.CLK(clknet_leaf_38_clk),
    .D(_01328_),
    .Q(\alu_shl[9] ));
 sky130_fd_sc_hd__dfxtp_1 _30832_ (.CLK(clknet_leaf_38_clk),
    .D(_01329_),
    .Q(\alu_shl[10] ));
 sky130_fd_sc_hd__dfxtp_1 _30833_ (.CLK(clknet_leaf_9_clk),
    .D(_01330_),
    .Q(\alu_shl[11] ));
 sky130_fd_sc_hd__dfxtp_1 _30834_ (.CLK(clknet_leaf_9_clk),
    .D(_01331_),
    .Q(\alu_shl[12] ));
 sky130_fd_sc_hd__dfxtp_1 _30835_ (.CLK(clknet_leaf_9_clk),
    .D(_01332_),
    .Q(\alu_shl[13] ));
 sky130_fd_sc_hd__dfxtp_1 _30836_ (.CLK(clknet_leaf_9_clk),
    .D(_01333_),
    .Q(\alu_shl[14] ));
 sky130_fd_sc_hd__dfxtp_1 _30837_ (.CLK(clknet_leaf_9_clk),
    .D(_01334_),
    .Q(\alu_shl[15] ));
 sky130_fd_sc_hd__dfxtp_2 _30838_ (.CLK(clknet_leaf_28_clk),
    .D(_01335_),
    .Q(\decoded_imm[31] ));
 sky130_fd_sc_hd__dfxtp_2 _30839_ (.CLK(clknet_leaf_27_clk),
    .D(_01336_),
    .Q(\decoded_imm[30] ));
 sky130_fd_sc_hd__dfxtp_2 _30840_ (.CLK(clknet_leaf_27_clk),
    .D(_01337_),
    .Q(\decoded_imm[29] ));
 sky130_fd_sc_hd__dfxtp_2 _30841_ (.CLK(clknet_leaf_27_clk),
    .D(_01338_),
    .Q(\decoded_imm[28] ));
 sky130_fd_sc_hd__dfxtp_2 _30842_ (.CLK(clknet_leaf_27_clk),
    .D(_01339_),
    .Q(\decoded_imm[27] ));
 sky130_fd_sc_hd__dfxtp_2 _30843_ (.CLK(clknet_leaf_27_clk),
    .D(_01340_),
    .Q(\decoded_imm[26] ));
 sky130_fd_sc_hd__dfxtp_2 _30844_ (.CLK(clknet_leaf_28_clk),
    .D(_01341_),
    .Q(\decoded_imm[25] ));
 sky130_fd_sc_hd__dfxtp_2 _30845_ (.CLK(clknet_leaf_28_clk),
    .D(_01342_),
    .Q(\decoded_imm[24] ));
 sky130_fd_sc_hd__dfxtp_1 _30846_ (.CLK(clknet_leaf_17_clk),
    .D(_01343_),
    .Q(\decoded_imm[23] ));
 sky130_fd_sc_hd__dfxtp_2 _30847_ (.CLK(clknet_leaf_27_clk),
    .D(_01344_),
    .Q(\decoded_imm[22] ));
 sky130_fd_sc_hd__dfxtp_2 _30848_ (.CLK(clknet_leaf_27_clk),
    .D(_01345_),
    .Q(\decoded_imm[21] ));
 sky130_fd_sc_hd__dfxtp_2 _30849_ (.CLK(clknet_leaf_27_clk),
    .D(_01346_),
    .Q(\decoded_imm[20] ));
 sky130_fd_sc_hd__dfxtp_2 _30850_ (.CLK(clknet_leaf_25_clk),
    .D(_01347_),
    .Q(\decoded_imm[19] ));
 sky130_fd_sc_hd__dfxtp_2 _30851_ (.CLK(clknet_leaf_25_clk),
    .D(_01348_),
    .Q(\decoded_imm[18] ));
 sky130_fd_sc_hd__dfxtp_1 _30852_ (.CLK(clknet_leaf_25_clk),
    .D(_01349_),
    .Q(\decoded_imm[17] ));
 sky130_fd_sc_hd__dfxtp_1 _30853_ (.CLK(clknet_leaf_25_clk),
    .D(_01350_),
    .Q(\decoded_imm[16] ));
 sky130_fd_sc_hd__dfxtp_1 _30854_ (.CLK(clknet_leaf_26_clk),
    .D(_01351_),
    .Q(\decoded_imm[15] ));
 sky130_fd_sc_hd__dfxtp_1 _30855_ (.CLK(clknet_leaf_26_clk),
    .D(_01352_),
    .Q(\decoded_imm[14] ));
 sky130_fd_sc_hd__dfxtp_1 _30856_ (.CLK(clknet_leaf_26_clk),
    .D(_01353_),
    .Q(\decoded_imm[13] ));
 sky130_fd_sc_hd__dfxtp_1 _30857_ (.CLK(clknet_leaf_26_clk),
    .D(_01354_),
    .Q(\decoded_imm[12] ));
 sky130_fd_sc_hd__dfxtp_2 _30858_ (.CLK(clknet_leaf_26_clk),
    .D(_01355_),
    .Q(\decoded_imm[11] ));
 sky130_fd_sc_hd__dfxtp_1 _30859_ (.CLK(clknet_leaf_26_clk),
    .D(_01356_),
    .Q(\decoded_imm[10] ));
 sky130_fd_sc_hd__dfxtp_2 _30860_ (.CLK(clknet_leaf_29_clk),
    .D(_01357_),
    .Q(\decoded_imm[9] ));
 sky130_fd_sc_hd__dfxtp_2 _30861_ (.CLK(clknet_leaf_25_clk),
    .D(_01358_),
    .Q(\decoded_imm[8] ));
 sky130_fd_sc_hd__dfxtp_1 _30862_ (.CLK(clknet_leaf_24_clk),
    .D(_01359_),
    .Q(\decoded_imm[7] ));
 sky130_fd_sc_hd__dfxtp_2 _30863_ (.CLK(clknet_leaf_29_clk),
    .D(_01360_),
    .Q(\decoded_imm[6] ));
 sky130_fd_sc_hd__dfxtp_1 _30864_ (.CLK(clknet_leaf_28_clk),
    .D(_01361_),
    .Q(\decoded_imm[5] ));
 sky130_fd_sc_hd__dfxtp_1 _30865_ (.CLK(clknet_leaf_28_clk),
    .D(_01362_),
    .Q(\decoded_imm[4] ));
 sky130_fd_sc_hd__dfxtp_2 _30866_ (.CLK(clknet_leaf_30_clk),
    .D(_01363_),
    .Q(\decoded_imm[3] ));
 sky130_fd_sc_hd__dfxtp_2 _30867_ (.CLK(clknet_leaf_31_clk),
    .D(_01364_),
    .Q(\decoded_imm[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30868_ (.CLK(clknet_leaf_33_clk),
    .D(_01365_),
    .Q(\decoded_imm[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30869_ (.CLK(clknet_leaf_89_clk),
    .D(_01366_),
    .Q(alu_wait));
 sky130_fd_sc_hd__dfxtp_1 _30870_ (.CLK(clknet_leaf_109_clk),
    .D(_01367_),
    .Q(\latched_rd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30871_ (.CLK(clknet_leaf_104_clk),
    .D(_01368_),
    .Q(\latched_rd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30872_ (.CLK(clknet_leaf_105_clk),
    .D(_01369_),
    .Q(\latched_rd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30873_ (.CLK(clknet_leaf_104_clk),
    .D(_01370_),
    .Q(\latched_rd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30874_ (.CLK(clknet_leaf_90_clk),
    .D(_01371_),
    .Q(\reg_next_pc[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30875_ (.CLK(clknet_leaf_173_clk),
    .D(_01372_),
    .Q(\cpuregs[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30876_ (.CLK(clknet_leaf_172_clk),
    .D(_01373_),
    .Q(\cpuregs[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30877_ (.CLK(clknet_leaf_172_clk),
    .D(_01374_),
    .Q(\cpuregs[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30878_ (.CLK(clknet_leaf_172_clk),
    .D(_01375_),
    .Q(\cpuregs[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30879_ (.CLK(clknet_leaf_173_clk),
    .D(_01376_),
    .Q(\cpuregs[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30880_ (.CLK(clknet_leaf_173_clk),
    .D(_01377_),
    .Q(\cpuregs[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30881_ (.CLK(clknet_leaf_180_clk),
    .D(_01378_),
    .Q(\cpuregs[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30882_ (.CLK(clknet_leaf_179_clk),
    .D(_01379_),
    .Q(\cpuregs[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30883_ (.CLK(clknet_leaf_170_clk),
    .D(_01380_),
    .Q(\cpuregs[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30884_ (.CLK(clknet_leaf_170_clk),
    .D(_01381_),
    .Q(\cpuregs[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30885_ (.CLK(clknet_leaf_179_clk),
    .D(_01382_),
    .Q(\cpuregs[19][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30886_ (.CLK(clknet_leaf_180_clk),
    .D(_01383_),
    .Q(\cpuregs[19][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30887_ (.CLK(clknet_leaf_101_clk),
    .D(_01384_),
    .Q(\cpuregs[19][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30888_ (.CLK(clknet_leaf_101_clk),
    .D(_01385_),
    .Q(\cpuregs[19][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30889_ (.CLK(clknet_leaf_99_clk),
    .D(_01386_),
    .Q(\cpuregs[19][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30890_ (.CLK(clknet_leaf_100_clk),
    .D(_01387_),
    .Q(\cpuregs[19][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30891_ (.CLK(clknet_leaf_103_clk),
    .D(_01388_),
    .Q(\cpuregs[19][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30892_ (.CLK(clknet_leaf_103_clk),
    .D(_01389_),
    .Q(\cpuregs[19][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30893_ (.CLK(clknet_leaf_160_clk),
    .D(_01390_),
    .Q(\cpuregs[19][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30894_ (.CLK(clknet_leaf_162_clk),
    .D(_01391_),
    .Q(\cpuregs[19][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30895_ (.CLK(clknet_leaf_163_clk),
    .D(_01392_),
    .Q(\cpuregs[19][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30896_ (.CLK(clknet_leaf_163_clk),
    .D(_01393_),
    .Q(\cpuregs[19][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30897_ (.CLK(clknet_leaf_163_clk),
    .D(_01394_),
    .Q(\cpuregs[19][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30898_ (.CLK(clknet_leaf_160_clk),
    .D(_01395_),
    .Q(\cpuregs[19][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30899_ (.CLK(clknet_leaf_120_clk),
    .D(_01396_),
    .Q(\cpuregs[19][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30900_ (.CLK(clknet_leaf_119_clk),
    .D(_01397_),
    .Q(\cpuregs[19][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30901_ (.CLK(clknet_leaf_115_clk),
    .D(_01398_),
    .Q(\cpuregs[19][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30902_ (.CLK(clknet_leaf_116_clk),
    .D(_01399_),
    .Q(\cpuregs[19][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30903_ (.CLK(clknet_leaf_121_clk),
    .D(_01400_),
    .Q(\cpuregs[19][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30904_ (.CLK(clknet_leaf_116_clk),
    .D(_01401_),
    .Q(\cpuregs[19][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30905_ (.CLK(clknet_leaf_121_clk),
    .D(_01402_),
    .Q(\cpuregs[19][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30906_ (.CLK(clknet_leaf_99_clk),
    .D(_01403_),
    .Q(\cpuregs[19][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30907_ (.CLK(clknet_leaf_105_clk),
    .D(_01404_),
    .Q(\latched_rd[4] ));
 sky130_fd_sc_hd__dfxtp_1 _30908_ (.CLK(clknet_leaf_91_clk),
    .D(_01405_),
    .Q(\decoded_rs1[4] ));
 sky130_fd_sc_hd__dfxtp_2 _30909_ (.CLK(clknet_leaf_34_clk),
    .D(_01406_),
    .Q(net119));
 sky130_fd_sc_hd__dfxtp_2 _30910_ (.CLK(clknet_leaf_34_clk),
    .D(_01407_),
    .Q(net122));
 sky130_fd_sc_hd__dfxtp_2 _30911_ (.CLK(clknet_leaf_34_clk),
    .D(_01408_),
    .Q(net123));
 sky130_fd_sc_hd__dfxtp_1 _30912_ (.CLK(clknet_leaf_49_clk),
    .D(_01409_),
    .Q(net124));
 sky130_fd_sc_hd__dfxtp_2 _30913_ (.CLK(clknet_leaf_36_clk),
    .D(_01410_),
    .Q(net125));
 sky130_fd_sc_hd__dfxtp_1 _30914_ (.CLK(clknet_leaf_12_clk),
    .D(_01411_),
    .Q(net126));
 sky130_fd_sc_hd__dfxtp_1 _30915_ (.CLK(clknet_leaf_36_clk),
    .D(_01412_),
    .Q(net127));
 sky130_fd_sc_hd__dfxtp_2 _30916_ (.CLK(clknet_leaf_36_clk),
    .D(_01413_),
    .Q(net128));
 sky130_fd_sc_hd__dfxtp_2 _30917_ (.CLK(clknet_leaf_20_clk),
    .D(_01414_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_1 _30918_ (.CLK(clknet_leaf_12_clk),
    .D(_01415_),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_2 _30919_ (.CLK(clknet_leaf_18_clk),
    .D(_01416_),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_2 _30920_ (.CLK(clknet_leaf_18_clk),
    .D(_01417_),
    .Q(net102));
 sky130_fd_sc_hd__dfxtp_2 _30921_ (.CLK(clknet_leaf_18_clk),
    .D(_01418_),
    .Q(net103));
 sky130_fd_sc_hd__dfxtp_2 _30922_ (.CLK(clknet_leaf_18_clk),
    .D(_01419_),
    .Q(net104));
 sky130_fd_sc_hd__dfxtp_2 _30923_ (.CLK(clknet_leaf_18_clk),
    .D(_01420_),
    .Q(net105));
 sky130_fd_sc_hd__dfxtp_2 _30924_ (.CLK(clknet_leaf_212_clk),
    .D(_01421_),
    .Q(net106));
 sky130_fd_sc_hd__dfxtp_2 _30925_ (.CLK(clknet_leaf_212_clk),
    .D(_01422_),
    .Q(net107));
 sky130_fd_sc_hd__dfxtp_2 _30926_ (.CLK(clknet_leaf_210_clk),
    .D(_01423_),
    .Q(net108));
 sky130_fd_sc_hd__dfxtp_2 _30927_ (.CLK(clknet_leaf_210_clk),
    .D(_01424_),
    .Q(net109));
 sky130_fd_sc_hd__dfxtp_2 _30928_ (.CLK(clknet_leaf_205_clk),
    .D(_01425_),
    .Q(net110));
 sky130_fd_sc_hd__dfxtp_2 _30929_ (.CLK(clknet_leaf_205_clk),
    .D(_01426_),
    .Q(net111));
 sky130_fd_sc_hd__dfxtp_2 _30930_ (.CLK(clknet_leaf_204_clk),
    .D(_01427_),
    .Q(net112));
 sky130_fd_sc_hd__dfxtp_2 _30931_ (.CLK(clknet_leaf_210_clk),
    .D(_01428_),
    .Q(net113));
 sky130_fd_sc_hd__dfxtp_2 _30932_ (.CLK(clknet_leaf_208_clk),
    .D(_01429_),
    .Q(net114));
 sky130_fd_sc_hd__dfxtp_2 _30933_ (.CLK(clknet_leaf_210_clk),
    .D(_01430_),
    .Q(net115));
 sky130_fd_sc_hd__dfxtp_2 _30934_ (.CLK(clknet_leaf_209_clk),
    .D(_01431_),
    .Q(net116));
 sky130_fd_sc_hd__dfxtp_2 _30935_ (.CLK(clknet_leaf_210_clk),
    .D(_01432_),
    .Q(net117));
 sky130_fd_sc_hd__dfxtp_2 _30936_ (.CLK(clknet_leaf_208_clk),
    .D(_01433_),
    .Q(net118));
 sky130_fd_sc_hd__dfxtp_2 _30937_ (.CLK(clknet_leaf_209_clk),
    .D(_01434_),
    .Q(net120));
 sky130_fd_sc_hd__dfxtp_2 _30938_ (.CLK(clknet_leaf_18_clk),
    .D(_01435_),
    .Q(net121));
 sky130_fd_sc_hd__dfxtp_1 _30939_ (.CLK(clknet_leaf_83_clk),
    .D(_00040_),
    .Q(\cpu_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _30940_ (.CLK(clknet_leaf_82_clk),
    .D(_00041_),
    .Q(\cpu_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _30941_ (.CLK(clknet_leaf_81_clk),
    .D(_00042_),
    .Q(\cpu_state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _30942_ (.CLK(clknet_leaf_97_clk),
    .D(_00043_),
    .Q(\cpu_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _30943_ (.CLK(clknet_leaf_82_clk),
    .D(_00044_),
    .Q(\cpu_state[4] ));
 sky130_fd_sc_hd__dfxtp_2 _30944_ (.CLK(clknet_leaf_85_clk),
    .D(_00045_),
    .Q(\cpu_state[5] ));
 sky130_fd_sc_hd__dfxtp_1 _30945_ (.CLK(clknet_leaf_82_clk),
    .D(_00046_),
    .Q(\cpu_state[6] ));
 sky130_fd_sc_hd__dfxtp_1 _30946_ (.CLK(clknet_leaf_158_clk),
    .D(_01436_),
    .Q(\cpuregs[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30947_ (.CLK(clknet_leaf_178_clk),
    .D(_01437_),
    .Q(\cpuregs[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30948_ (.CLK(clknet_leaf_177_clk),
    .D(_01438_),
    .Q(\cpuregs[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30949_ (.CLK(clknet_leaf_186_clk),
    .D(_01439_),
    .Q(\cpuregs[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30950_ (.CLK(clknet_leaf_178_clk),
    .D(_01440_),
    .Q(\cpuregs[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30951_ (.CLK(clknet_leaf_169_clk),
    .D(_01441_),
    .Q(\cpuregs[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30952_ (.CLK(clknet_leaf_188_clk),
    .D(_01442_),
    .Q(\cpuregs[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30953_ (.CLK(clknet_leaf_191_clk),
    .D(_01443_),
    .Q(\cpuregs[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30954_ (.CLK(clknet_leaf_156_clk),
    .D(_01444_),
    .Q(\cpuregs[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30955_ (.CLK(clknet_leaf_154_clk),
    .D(_01445_),
    .Q(\cpuregs[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30956_ (.CLK(clknet_leaf_191_clk),
    .D(_01446_),
    .Q(\cpuregs[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30957_ (.CLK(clknet_leaf_189_clk),
    .D(_01447_),
    .Q(\cpuregs[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30958_ (.CLK(clknet_leaf_137_clk),
    .D(_01448_),
    .Q(\cpuregs[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30959_ (.CLK(clknet_leaf_140_clk),
    .D(_01449_),
    .Q(\cpuregs[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30960_ (.CLK(clknet_leaf_164_clk),
    .D(_01450_),
    .Q(\cpuregs[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30961_ (.CLK(clknet_leaf_142_clk),
    .D(_01451_),
    .Q(\cpuregs[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30962_ (.CLK(clknet_leaf_137_clk),
    .D(_01452_),
    .Q(\cpuregs[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30963_ (.CLK(clknet_leaf_124_clk),
    .D(_01453_),
    .Q(\cpuregs[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30964_ (.CLK(clknet_leaf_143_clk),
    .D(_01454_),
    .Q(\cpuregs[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30965_ (.CLK(clknet_leaf_149_clk),
    .D(_01455_),
    .Q(\cpuregs[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30966_ (.CLK(clknet_leaf_149_clk),
    .D(_01456_),
    .Q(\cpuregs[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30967_ (.CLK(clknet_leaf_148_clk),
    .D(_01457_),
    .Q(\cpuregs[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _30968_ (.CLK(clknet_leaf_147_clk),
    .D(_01458_),
    .Q(\cpuregs[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _30969_ (.CLK(clknet_leaf_161_clk),
    .D(_01459_),
    .Q(\cpuregs[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _30970_ (.CLK(clknet_leaf_132_clk),
    .D(_01460_),
    .Q(\cpuregs[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _30971_ (.CLK(clknet_leaf_132_clk),
    .D(_01461_),
    .Q(\cpuregs[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _30972_ (.CLK(clknet_leaf_121_clk),
    .D(_01462_),
    .Q(\cpuregs[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _30973_ (.CLK(clknet_leaf_118_clk),
    .D(_01463_),
    .Q(\cpuregs[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _30974_ (.CLK(clknet_leaf_126_clk),
    .D(_01464_),
    .Q(\cpuregs[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _30975_ (.CLK(clknet_leaf_118_clk),
    .D(_01465_),
    .Q(\cpuregs[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _30976_ (.CLK(clknet_leaf_138_clk),
    .D(_01466_),
    .Q(\cpuregs[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _30977_ (.CLK(clknet_leaf_142_clk),
    .D(_01467_),
    .Q(\cpuregs[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 _30978_ (.CLK(clknet_leaf_159_clk),
    .D(_01468_),
    .Q(\cpuregs[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _30979_ (.CLK(clknet_leaf_172_clk),
    .D(_01469_),
    .Q(\cpuregs[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _30980_ (.CLK(clknet_leaf_172_clk),
    .D(_01470_),
    .Q(\cpuregs[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _30981_ (.CLK(clknet_leaf_168_clk),
    .D(_01471_),
    .Q(\cpuregs[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _30982_ (.CLK(clknet_leaf_170_clk),
    .D(_01472_),
    .Q(\cpuregs[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _30983_ (.CLK(clknet_leaf_168_clk),
    .D(_01473_),
    .Q(\cpuregs[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _30984_ (.CLK(clknet_leaf_185_clk),
    .D(_01474_),
    .Q(\cpuregs[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _30985_ (.CLK(clknet_leaf_193_clk),
    .D(_01475_),
    .Q(\cpuregs[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _30986_ (.CLK(clknet_leaf_192_clk),
    .D(_01476_),
    .Q(\cpuregs[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _30987_ (.CLK(clknet_leaf_192_clk),
    .D(_01477_),
    .Q(\cpuregs[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _30988_ (.CLK(clknet_leaf_190_clk),
    .D(_01478_),
    .Q(\cpuregs[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _30989_ (.CLK(clknet_leaf_188_clk),
    .D(_01479_),
    .Q(\cpuregs[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _30990_ (.CLK(clknet_leaf_139_clk),
    .D(_01480_),
    .Q(\cpuregs[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _30991_ (.CLK(clknet_leaf_100_clk),
    .D(_01481_),
    .Q(\cpuregs[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _30992_ (.CLK(clknet_leaf_100_clk),
    .D(_01482_),
    .Q(\cpuregs[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _30993_ (.CLK(clknet_leaf_164_clk),
    .D(_01483_),
    .Q(\cpuregs[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _30994_ (.CLK(clknet_leaf_124_clk),
    .D(_01484_),
    .Q(\cpuregs[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _30995_ (.CLK(clknet_leaf_121_clk),
    .D(_01485_),
    .Q(\cpuregs[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _30996_ (.CLK(clknet_leaf_143_clk),
    .D(_01486_),
    .Q(\cpuregs[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _30997_ (.CLK(clknet_leaf_162_clk),
    .D(_01487_),
    .Q(\cpuregs[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _30998_ (.CLK(clknet_leaf_162_clk),
    .D(_01488_),
    .Q(\cpuregs[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _30999_ (.CLK(clknet_leaf_162_clk),
    .D(_01489_),
    .Q(\cpuregs[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _31000_ (.CLK(clknet_leaf_143_clk),
    .D(_01490_),
    .Q(\cpuregs[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _31001_ (.CLK(clknet_leaf_162_clk),
    .D(_01491_),
    .Q(\cpuregs[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _31002_ (.CLK(clknet_leaf_124_clk),
    .D(_01492_),
    .Q(\cpuregs[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _31003_ (.CLK(clknet_leaf_125_clk),
    .D(_01493_),
    .Q(\cpuregs[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _31004_ (.CLK(clknet_leaf_116_clk),
    .D(_01494_),
    .Q(\cpuregs[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _31005_ (.CLK(clknet_leaf_120_clk),
    .D(_01495_),
    .Q(\cpuregs[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _31006_ (.CLK(clknet_leaf_125_clk),
    .D(_01496_),
    .Q(\cpuregs[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _31007_ (.CLK(clknet_leaf_116_clk),
    .D(_01497_),
    .Q(\cpuregs[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _31008_ (.CLK(clknet_leaf_134_clk),
    .D(_01498_),
    .Q(\cpuregs[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _31009_ (.CLK(clknet_leaf_141_clk),
    .D(_01499_),
    .Q(\cpuregs[1][31] ));
 sky130_fd_sc_hd__conb_1 picorv32a_375 (.LO(net375));
 sky130_fd_sc_hd__conb_1 picorv32a_376 (.LO(net376));
 sky130_fd_sc_hd__conb_1 picorv32a_377 (.LO(net377));
 sky130_fd_sc_hd__conb_1 picorv32a_378 (.LO(net378));
 sky130_fd_sc_hd__conb_1 picorv32a_379 (.LO(net379));
 sky130_fd_sc_hd__conb_1 picorv32a_380 (.LO(net380));
 sky130_fd_sc_hd__conb_1 picorv32a_381 (.LO(net381));
 sky130_fd_sc_hd__conb_1 picorv32a_382 (.LO(net382));
 sky130_fd_sc_hd__conb_1 picorv32a_383 (.LO(net383));
 sky130_fd_sc_hd__conb_1 picorv32a_384 (.LO(net384));
 sky130_fd_sc_hd__conb_1 picorv32a_385 (.LO(net385));
 sky130_fd_sc_hd__conb_1 picorv32a_386 (.LO(net386));
 sky130_fd_sc_hd__conb_1 picorv32a_387 (.LO(net387));
 sky130_fd_sc_hd__conb_1 picorv32a_388 (.LO(net388));
 sky130_fd_sc_hd__conb_1 picorv32a_389 (.LO(net389));
 sky130_fd_sc_hd__conb_1 picorv32a_390 (.LO(net390));
 sky130_fd_sc_hd__conb_1 picorv32a_391 (.LO(net391));
 sky130_fd_sc_hd__conb_1 picorv32a_392 (.LO(net392));
 sky130_fd_sc_hd__conb_1 picorv32a_393 (.LO(net393));
 sky130_fd_sc_hd__conb_1 picorv32a_394 (.LO(net394));
 sky130_fd_sc_hd__conb_1 picorv32a_395 (.LO(net395));
 sky130_fd_sc_hd__conb_1 picorv32a_396 (.LO(net396));
 sky130_fd_sc_hd__conb_1 picorv32a_397 (.LO(net397));
 sky130_fd_sc_hd__conb_1 picorv32a_398 (.LO(net398));
 sky130_fd_sc_hd__conb_1 picorv32a_399 (.LO(net399));
 sky130_fd_sc_hd__conb_1 picorv32a_400 (.LO(net400));
 sky130_fd_sc_hd__conb_1 picorv32a_401 (.LO(net401));
 sky130_fd_sc_hd__conb_1 picorv32a_402 (.LO(net402));
 sky130_fd_sc_hd__conb_1 picorv32a_403 (.LO(net403));
 sky130_fd_sc_hd__conb_1 picorv32a_404 (.LO(net404));
 sky130_fd_sc_hd__conb_1 picorv32a_405 (.LO(net405));
 sky130_fd_sc_hd__conb_1 picorv32a_406 (.LO(net406));
 sky130_fd_sc_hd__conb_1 picorv32a_407 (.LO(net407));
 sky130_fd_sc_hd__conb_1 picorv32a_408 (.LO(net408));
 sky130_fd_sc_hd__conb_1 picorv32a_409 (.LO(net409));
 sky130_fd_sc_hd__conb_1 picorv32a_410 (.LO(net410));
 sky130_fd_sc_hd__conb_1 picorv32a_411 (.LO(net411));
 sky130_fd_sc_hd__conb_1 picorv32a_412 (.LO(net412));
 sky130_fd_sc_hd__conb_1 picorv32a_413 (.LO(net413));
 sky130_fd_sc_hd__conb_1 picorv32a_414 (.LO(net414));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__buf_1 _31051_ (.A(net161),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_1 _31052_ (.A(net172),
    .X(net310));
 sky130_fd_sc_hd__buf_2 _31053_ (.A(net183),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_2 _31054_ (.A(net186),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_2 _31055_ (.A(net187),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_4 _31056_ (.A(net188),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_4 _31057_ (.A(net189),
    .X(net327));
 sky130_fd_sc_hd__buf_1 _31058_ (.A(net190),
    .X(net328));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Right_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Right_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Right_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Right_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Right_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Right_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Right_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Right_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Right_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Right_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Right_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Right_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Right_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Right_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Right_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Right_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Right_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Right_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Right_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Right_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Right_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Right_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Right_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Right_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Right_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Right_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Right_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Right_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Right_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Right_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Right_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Right_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Right_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_Right_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_Right_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_Right_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_Right_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_Right_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_Right_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_Right_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_Right_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_Right_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_Right_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_Right_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_Right_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_Right_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_Right_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_Right_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_Right_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_Right_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_Right_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_Right_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_Right_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_Right_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_Right_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_Right_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_Right_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_Right_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_Right_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_Right_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_Right_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_Right_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_Right_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_Right_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_228_Right_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_229_Right_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_230_Right_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_231_Right_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_232_Right_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_233_Right_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_234_Right_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_235_Right_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_236_Right_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_237_Right_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_238_Right_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_239_Right_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_240_Right_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_241_Right_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_242_Right_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_243_Right_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_244_Right_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_245_Right_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_246_Right_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_247_Right_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_248_Right_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_249_Right_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_333 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_334 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_335 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_336 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_337 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_338 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_339 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_340 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_341 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_342 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_343 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_344 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_345 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_346 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_347 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_348 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_349 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_350 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_351 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_352 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_353 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_354 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_355 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_356 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_357 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_358 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_359 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_360 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_361 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_362 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_363 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_364 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_365 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_366 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_367 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_368 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_369 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_370 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_371 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_372 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_373 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_374 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_375 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_376 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_377 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_378 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_379 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_380 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_381 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_382 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_383 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_384 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_385 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_386 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_387 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_388 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_389 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_390 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_391 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_392 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_393 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_394 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_395 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_396 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_397 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_398 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_399 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_400 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_401 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_402 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_403 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_404 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Left_405 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Left_406 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Left_407 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Left_408 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Left_409 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Left_410 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Left_411 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Left_412 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Left_413 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Left_414 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Left_415 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Left_416 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Left_417 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Left_418 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Left_419 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Left_420 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Left_421 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Left_422 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Left_423 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Left_424 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Left_425 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Left_426 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Left_427 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Left_428 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Left_429 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Left_430 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Left_431 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Left_432 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Left_433 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Left_434 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Left_435 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Left_436 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Left_437 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Left_438 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Left_439 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Left_440 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Left_441 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Left_442 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Left_443 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Left_444 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Left_445 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Left_446 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_Left_447 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_Left_448 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_Left_449 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_Left_450 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_Left_451 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_Left_452 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_Left_453 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_Left_454 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_Left_455 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_Left_456 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_Left_457 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_Left_458 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_Left_459 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_Left_460 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_Left_461 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_Left_462 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_Left_463 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_Left_464 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_Left_465 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_Left_466 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_Left_467 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_Left_468 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_Left_469 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_Left_470 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_Left_471 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_Left_472 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_Left_473 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_Left_474 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_Left_475 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_Left_476 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_Left_477 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_228_Left_478 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_229_Left_479 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_230_Left_480 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_231_Left_481 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_232_Left_482 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_233_Left_483 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_234_Left_484 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_235_Left_485 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_236_Left_486 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_237_Left_487 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_238_Left_488 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_239_Left_489 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_240_Left_490 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_241_Left_491 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_242_Left_492 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_243_Left_493 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_244_Left_494 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_245_Left_495 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_246_Left_496 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_247_Left_497 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_248_Left_498 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_249_Left_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_7051 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(irq[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(irq[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(irq[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(irq[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(irq[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(irq[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(irq[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(irq[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(irq[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(irq[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(irq[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(irq[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(irq[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(irq[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(irq[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(irq[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(irq[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(irq[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(irq[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(irq[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(irq[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(irq[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(irq[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(irq[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(irq[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(irq[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(irq[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(irq[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(irq[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(irq[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(irq[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(irq[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_2 input33 (.A(mem_rdata[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(mem_rdata[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(mem_rdata[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(mem_rdata[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_2 input37 (.A(mem_rdata[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(mem_rdata[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_2 input39 (.A(mem_rdata[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(mem_rdata[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(mem_rdata[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(mem_rdata[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(mem_rdata[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(mem_rdata[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_2 input45 (.A(mem_rdata[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_2 input46 (.A(mem_rdata[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_2 input47 (.A(mem_rdata[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(mem_rdata[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_2 input49 (.A(mem_rdata[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_2 input50 (.A(mem_rdata[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_2 input51 (.A(mem_rdata[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_2 input52 (.A(mem_rdata[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(mem_rdata[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_2 input54 (.A(mem_rdata[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(mem_rdata[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_2 input56 (.A(mem_rdata[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(mem_rdata[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(mem_rdata[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(mem_rdata[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(mem_rdata[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(mem_rdata[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(mem_rdata[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_2 input63 (.A(mem_rdata[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 input64 (.A(mem_rdata[9]),
    .X(net64));
 sky130_fd_sc_hd__dlymetal6s2s_1 input65 (.A(mem_ready),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(resetn),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net67),
    .X(eoi[0]));
 sky130_fd_sc_hd__clkbuf_4 output68 (.A(net68),
    .X(eoi[10]));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net69),
    .X(eoi[11]));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net70),
    .X(eoi[12]));
 sky130_fd_sc_hd__clkbuf_4 output71 (.A(net71),
    .X(eoi[13]));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net72),
    .X(eoi[14]));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net73),
    .X(eoi[15]));
 sky130_fd_sc_hd__clkbuf_4 output74 (.A(net74),
    .X(eoi[16]));
 sky130_fd_sc_hd__clkbuf_4 output75 (.A(net75),
    .X(eoi[17]));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net76),
    .X(eoi[18]));
 sky130_fd_sc_hd__clkbuf_4 output77 (.A(net77),
    .X(eoi[19]));
 sky130_fd_sc_hd__clkbuf_4 output78 (.A(net78),
    .X(eoi[1]));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net79),
    .X(eoi[20]));
 sky130_fd_sc_hd__clkbuf_4 output80 (.A(net80),
    .X(eoi[21]));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net81),
    .X(eoi[22]));
 sky130_fd_sc_hd__clkbuf_4 output82 (.A(net82),
    .X(eoi[23]));
 sky130_fd_sc_hd__clkbuf_4 output83 (.A(net83),
    .X(eoi[24]));
 sky130_fd_sc_hd__clkbuf_4 output84 (.A(net84),
    .X(eoi[25]));
 sky130_fd_sc_hd__clkbuf_4 output85 (.A(net85),
    .X(eoi[26]));
 sky130_fd_sc_hd__clkbuf_4 output86 (.A(net86),
    .X(eoi[27]));
 sky130_fd_sc_hd__clkbuf_4 output87 (.A(net87),
    .X(eoi[28]));
 sky130_fd_sc_hd__clkbuf_4 output88 (.A(net88),
    .X(eoi[29]));
 sky130_fd_sc_hd__clkbuf_4 output89 (.A(net89),
    .X(eoi[2]));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net90),
    .X(eoi[30]));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net91),
    .X(eoi[31]));
 sky130_fd_sc_hd__clkbuf_4 output92 (.A(net92),
    .X(eoi[3]));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net93),
    .X(eoi[4]));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net94),
    .X(eoi[5]));
 sky130_fd_sc_hd__clkbuf_4 output95 (.A(net95),
    .X(eoi[6]));
 sky130_fd_sc_hd__clkbuf_4 output96 (.A(net96),
    .X(eoi[7]));
 sky130_fd_sc_hd__clkbuf_4 output97 (.A(net97),
    .X(eoi[8]));
 sky130_fd_sc_hd__clkbuf_4 output98 (.A(net98),
    .X(eoi[9]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(mem_addr[10]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(mem_addr[11]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(mem_addr[12]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(mem_addr[13]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(mem_addr[14]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(mem_addr[15]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(mem_addr[16]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(mem_addr[17]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(mem_addr[18]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(mem_addr[19]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(mem_addr[20]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(mem_addr[21]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(mem_addr[22]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(mem_addr[23]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(mem_addr[24]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(mem_addr[25]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(mem_addr[26]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(mem_addr[27]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(mem_addr[28]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(mem_addr[29]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(mem_addr[2]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(mem_addr[30]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(mem_addr[31]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(mem_addr[3]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(mem_addr[4]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(mem_addr[5]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(mem_addr[6]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(mem_addr[7]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(mem_addr[8]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(mem_addr[9]));
 sky130_fd_sc_hd__clkbuf_4 output129 (.A(net129),
    .X(mem_instr));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(mem_la_addr[10]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(mem_la_addr[11]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(mem_la_addr[12]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(mem_la_addr[13]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(mem_la_addr[14]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(mem_la_addr[15]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(mem_la_addr[16]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net137),
    .X(mem_la_addr[17]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(mem_la_addr[18]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(mem_la_addr[19]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(mem_la_addr[20]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(mem_la_addr[21]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(mem_la_addr[22]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net143),
    .X(mem_la_addr[23]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net144),
    .X(mem_la_addr[24]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net145),
    .X(mem_la_addr[25]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(mem_la_addr[26]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net147),
    .X(mem_la_addr[27]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net148),
    .X(mem_la_addr[28]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net149),
    .X(mem_la_addr[29]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net150),
    .X(mem_la_addr[2]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net151),
    .X(mem_la_addr[30]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net152),
    .X(mem_la_addr[31]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net153),
    .X(mem_la_addr[3]));
 sky130_fd_sc_hd__clkbuf_4 output154 (.A(net154),
    .X(mem_la_addr[4]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(mem_la_addr[5]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(mem_la_addr[6]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(mem_la_addr[7]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(mem_la_addr[8]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(mem_la_addr[9]));
 sky130_fd_sc_hd__clkbuf_4 output160 (.A(net160),
    .X(mem_la_read));
 sky130_fd_sc_hd__buf_2 output161 (.A(net161),
    .X(mem_la_wdata[0]));
 sky130_fd_sc_hd__buf_2 output162 (.A(net162),
    .X(mem_la_wdata[10]));
 sky130_fd_sc_hd__clkbuf_4 output163 (.A(net163),
    .X(mem_la_wdata[11]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net164),
    .X(mem_la_wdata[12]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net165),
    .X(mem_la_wdata[13]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(mem_la_wdata[14]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(mem_la_wdata[15]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(mem_la_wdata[16]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net169),
    .X(mem_la_wdata[17]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net170),
    .X(mem_la_wdata[18]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net171),
    .X(mem_la_wdata[19]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(mem_la_wdata[1]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net173),
    .X(mem_la_wdata[20]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net174),
    .X(mem_la_wdata[21]));
 sky130_fd_sc_hd__buf_2 output175 (.A(net175),
    .X(mem_la_wdata[22]));
 sky130_fd_sc_hd__buf_2 output176 (.A(net176),
    .X(mem_la_wdata[23]));
 sky130_fd_sc_hd__buf_2 output177 (.A(net177),
    .X(mem_la_wdata[24]));
 sky130_fd_sc_hd__buf_2 output178 (.A(net178),
    .X(mem_la_wdata[25]));
 sky130_fd_sc_hd__buf_2 output179 (.A(net179),
    .X(mem_la_wdata[26]));
 sky130_fd_sc_hd__buf_2 output180 (.A(net180),
    .X(mem_la_wdata[27]));
 sky130_fd_sc_hd__buf_2 output181 (.A(net181),
    .X(mem_la_wdata[28]));
 sky130_fd_sc_hd__buf_2 output182 (.A(net182),
    .X(mem_la_wdata[29]));
 sky130_fd_sc_hd__buf_2 output183 (.A(net183),
    .X(mem_la_wdata[2]));
 sky130_fd_sc_hd__buf_2 output184 (.A(net184),
    .X(mem_la_wdata[30]));
 sky130_fd_sc_hd__buf_2 output185 (.A(net185),
    .X(mem_la_wdata[31]));
 sky130_fd_sc_hd__buf_2 output186 (.A(net186),
    .X(mem_la_wdata[3]));
 sky130_fd_sc_hd__buf_2 output187 (.A(net187),
    .X(mem_la_wdata[4]));
 sky130_fd_sc_hd__buf_2 output188 (.A(net188),
    .X(mem_la_wdata[5]));
 sky130_fd_sc_hd__buf_2 output189 (.A(net189),
    .X(mem_la_wdata[6]));
 sky130_fd_sc_hd__buf_2 output190 (.A(net190),
    .X(mem_la_wdata[7]));
 sky130_fd_sc_hd__buf_2 output191 (.A(net191),
    .X(mem_la_wdata[8]));
 sky130_fd_sc_hd__buf_2 output192 (.A(net192),
    .X(mem_la_wdata[9]));
 sky130_fd_sc_hd__clkbuf_4 output193 (.A(net193),
    .X(mem_la_write));
 sky130_fd_sc_hd__buf_2 output194 (.A(net194),
    .X(mem_la_wstrb[0]));
 sky130_fd_sc_hd__clkbuf_4 output195 (.A(net195),
    .X(mem_la_wstrb[1]));
 sky130_fd_sc_hd__clkbuf_4 output196 (.A(net196),
    .X(mem_la_wstrb[2]));
 sky130_fd_sc_hd__clkbuf_4 output197 (.A(net197),
    .X(mem_la_wstrb[3]));
 sky130_fd_sc_hd__clkbuf_4 output198 (.A(net198),
    .X(mem_valid));
 sky130_fd_sc_hd__clkbuf_4 output199 (.A(net199),
    .X(mem_wdata[0]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net200),
    .X(mem_wdata[10]));
 sky130_fd_sc_hd__buf_2 output201 (.A(net201),
    .X(mem_wdata[11]));
 sky130_fd_sc_hd__buf_2 output202 (.A(net202),
    .X(mem_wdata[12]));
 sky130_fd_sc_hd__buf_2 output203 (.A(net203),
    .X(mem_wdata[13]));
 sky130_fd_sc_hd__buf_2 output204 (.A(net204),
    .X(mem_wdata[14]));
 sky130_fd_sc_hd__buf_2 output205 (.A(net205),
    .X(mem_wdata[15]));
 sky130_fd_sc_hd__buf_2 output206 (.A(net206),
    .X(mem_wdata[16]));
 sky130_fd_sc_hd__buf_2 output207 (.A(net207),
    .X(mem_wdata[17]));
 sky130_fd_sc_hd__buf_2 output208 (.A(net208),
    .X(mem_wdata[18]));
 sky130_fd_sc_hd__buf_2 output209 (.A(net209),
    .X(mem_wdata[19]));
 sky130_fd_sc_hd__clkbuf_4 output210 (.A(net210),
    .X(mem_wdata[1]));
 sky130_fd_sc_hd__buf_2 output211 (.A(net211),
    .X(mem_wdata[20]));
 sky130_fd_sc_hd__buf_2 output212 (.A(net212),
    .X(mem_wdata[21]));
 sky130_fd_sc_hd__buf_2 output213 (.A(net213),
    .X(mem_wdata[22]));
 sky130_fd_sc_hd__buf_2 output214 (.A(net214),
    .X(mem_wdata[23]));
 sky130_fd_sc_hd__buf_2 output215 (.A(net215),
    .X(mem_wdata[24]));
 sky130_fd_sc_hd__clkbuf_4 output216 (.A(net216),
    .X(mem_wdata[25]));
 sky130_fd_sc_hd__buf_2 output217 (.A(net217),
    .X(mem_wdata[26]));
 sky130_fd_sc_hd__buf_2 output218 (.A(net218),
    .X(mem_wdata[27]));
 sky130_fd_sc_hd__buf_2 output219 (.A(net219),
    .X(mem_wdata[28]));
 sky130_fd_sc_hd__buf_2 output220 (.A(net220),
    .X(mem_wdata[29]));
 sky130_fd_sc_hd__buf_2 output221 (.A(net221),
    .X(mem_wdata[2]));
 sky130_fd_sc_hd__buf_2 output222 (.A(net222),
    .X(mem_wdata[30]));
 sky130_fd_sc_hd__clkbuf_4 output223 (.A(net223),
    .X(mem_wdata[31]));
 sky130_fd_sc_hd__buf_2 output224 (.A(net224),
    .X(mem_wdata[3]));
 sky130_fd_sc_hd__buf_2 output225 (.A(net225),
    .X(mem_wdata[4]));
 sky130_fd_sc_hd__buf_2 output226 (.A(net226),
    .X(mem_wdata[5]));
 sky130_fd_sc_hd__buf_2 output227 (.A(net227),
    .X(mem_wdata[6]));
 sky130_fd_sc_hd__buf_2 output228 (.A(net228),
    .X(mem_wdata[7]));
 sky130_fd_sc_hd__buf_2 output229 (.A(net229),
    .X(mem_wdata[8]));
 sky130_fd_sc_hd__buf_2 output230 (.A(net230),
    .X(mem_wdata[9]));
 sky130_fd_sc_hd__clkbuf_4 output231 (.A(net231),
    .X(mem_wstrb[0]));
 sky130_fd_sc_hd__clkbuf_4 output232 (.A(net232),
    .X(mem_wstrb[1]));
 sky130_fd_sc_hd__clkbuf_4 output233 (.A(net233),
    .X(mem_wstrb[2]));
 sky130_fd_sc_hd__clkbuf_4 output234 (.A(net234),
    .X(mem_wstrb[3]));
 sky130_fd_sc_hd__clkbuf_4 output235 (.A(net235),
    .X(pcpi_insn[0]));
 sky130_fd_sc_hd__clkbuf_4 output236 (.A(net236),
    .X(pcpi_insn[10]));
 sky130_fd_sc_hd__clkbuf_4 output237 (.A(net237),
    .X(pcpi_insn[11]));
 sky130_fd_sc_hd__buf_2 output238 (.A(net238),
    .X(pcpi_insn[12]));
 sky130_fd_sc_hd__buf_2 output239 (.A(net239),
    .X(pcpi_insn[13]));
 sky130_fd_sc_hd__clkbuf_4 output240 (.A(net240),
    .X(pcpi_insn[14]));
 sky130_fd_sc_hd__clkbuf_4 output241 (.A(net241),
    .X(pcpi_insn[15]));
 sky130_fd_sc_hd__clkbuf_4 output242 (.A(net242),
    .X(pcpi_insn[16]));
 sky130_fd_sc_hd__clkbuf_4 output243 (.A(net243),
    .X(pcpi_insn[17]));
 sky130_fd_sc_hd__clkbuf_4 output244 (.A(net244),
    .X(pcpi_insn[18]));
 sky130_fd_sc_hd__clkbuf_4 output245 (.A(net245),
    .X(pcpi_insn[19]));
 sky130_fd_sc_hd__clkbuf_4 output246 (.A(net246),
    .X(pcpi_insn[1]));
 sky130_fd_sc_hd__clkbuf_4 output247 (.A(net247),
    .X(pcpi_insn[20]));
 sky130_fd_sc_hd__clkbuf_4 output248 (.A(net248),
    .X(pcpi_insn[21]));
 sky130_fd_sc_hd__clkbuf_4 output249 (.A(net249),
    .X(pcpi_insn[22]));
 sky130_fd_sc_hd__clkbuf_4 output250 (.A(net250),
    .X(pcpi_insn[23]));
 sky130_fd_sc_hd__buf_2 output251 (.A(net251),
    .X(pcpi_insn[24]));
 sky130_fd_sc_hd__clkbuf_4 output252 (.A(net252),
    .X(pcpi_insn[25]));
 sky130_fd_sc_hd__clkbuf_4 output253 (.A(net253),
    .X(pcpi_insn[26]));
 sky130_fd_sc_hd__clkbuf_4 output254 (.A(net254),
    .X(pcpi_insn[27]));
 sky130_fd_sc_hd__clkbuf_4 output255 (.A(net255),
    .X(pcpi_insn[28]));
 sky130_fd_sc_hd__buf_2 output256 (.A(net256),
    .X(pcpi_insn[29]));
 sky130_fd_sc_hd__clkbuf_4 output257 (.A(net257),
    .X(pcpi_insn[2]));
 sky130_fd_sc_hd__clkbuf_4 output258 (.A(net258),
    .X(pcpi_insn[30]));
 sky130_fd_sc_hd__buf_2 output259 (.A(net259),
    .X(pcpi_insn[31]));
 sky130_fd_sc_hd__clkbuf_4 output260 (.A(net260),
    .X(pcpi_insn[3]));
 sky130_fd_sc_hd__clkbuf_4 output261 (.A(net261),
    .X(pcpi_insn[4]));
 sky130_fd_sc_hd__clkbuf_4 output262 (.A(net262),
    .X(pcpi_insn[5]));
 sky130_fd_sc_hd__clkbuf_4 output263 (.A(net263),
    .X(pcpi_insn[6]));
 sky130_fd_sc_hd__clkbuf_4 output264 (.A(net264),
    .X(pcpi_insn[7]));
 sky130_fd_sc_hd__clkbuf_4 output265 (.A(net265),
    .X(pcpi_insn[8]));
 sky130_fd_sc_hd__clkbuf_4 output266 (.A(net266),
    .X(pcpi_insn[9]));
 sky130_fd_sc_hd__buf_2 output267 (.A(net267),
    .X(pcpi_rs1[0]));
 sky130_fd_sc_hd__buf_2 output268 (.A(net268),
    .X(pcpi_rs1[10]));
 sky130_fd_sc_hd__buf_2 output269 (.A(net269),
    .X(pcpi_rs1[11]));
 sky130_fd_sc_hd__buf_2 output270 (.A(net270),
    .X(pcpi_rs1[12]));
 sky130_fd_sc_hd__buf_2 output271 (.A(net271),
    .X(pcpi_rs1[13]));
 sky130_fd_sc_hd__buf_2 output272 (.A(net272),
    .X(pcpi_rs1[14]));
 sky130_fd_sc_hd__buf_2 output273 (.A(net273),
    .X(pcpi_rs1[15]));
 sky130_fd_sc_hd__buf_2 output274 (.A(net274),
    .X(pcpi_rs1[16]));
 sky130_fd_sc_hd__buf_2 output275 (.A(net275),
    .X(pcpi_rs1[17]));
 sky130_fd_sc_hd__buf_2 output276 (.A(net276),
    .X(pcpi_rs1[18]));
 sky130_fd_sc_hd__buf_2 output277 (.A(net277),
    .X(pcpi_rs1[19]));
 sky130_fd_sc_hd__buf_2 output278 (.A(net278),
    .X(pcpi_rs1[1]));
 sky130_fd_sc_hd__buf_2 output279 (.A(net279),
    .X(pcpi_rs1[20]));
 sky130_fd_sc_hd__buf_2 output280 (.A(net280),
    .X(pcpi_rs1[21]));
 sky130_fd_sc_hd__buf_2 output281 (.A(net281),
    .X(pcpi_rs1[22]));
 sky130_fd_sc_hd__buf_2 output282 (.A(net282),
    .X(pcpi_rs1[23]));
 sky130_fd_sc_hd__buf_2 output283 (.A(net283),
    .X(pcpi_rs1[24]));
 sky130_fd_sc_hd__buf_2 output284 (.A(net284),
    .X(pcpi_rs1[25]));
 sky130_fd_sc_hd__buf_2 output285 (.A(net285),
    .X(pcpi_rs1[26]));
 sky130_fd_sc_hd__buf_2 output286 (.A(net286),
    .X(pcpi_rs1[27]));
 sky130_fd_sc_hd__buf_2 output287 (.A(net287),
    .X(pcpi_rs1[28]));
 sky130_fd_sc_hd__buf_2 output288 (.A(net288),
    .X(pcpi_rs1[29]));
 sky130_fd_sc_hd__buf_2 output289 (.A(net289),
    .X(pcpi_rs1[2]));
 sky130_fd_sc_hd__buf_2 output290 (.A(net290),
    .X(pcpi_rs1[30]));
 sky130_fd_sc_hd__buf_2 output291 (.A(net291),
    .X(pcpi_rs1[31]));
 sky130_fd_sc_hd__buf_2 output292 (.A(net292),
    .X(pcpi_rs1[3]));
 sky130_fd_sc_hd__buf_2 output293 (.A(net293),
    .X(pcpi_rs1[4]));
 sky130_fd_sc_hd__buf_2 output294 (.A(net294),
    .X(pcpi_rs1[5]));
 sky130_fd_sc_hd__buf_2 output295 (.A(net295),
    .X(pcpi_rs1[6]));
 sky130_fd_sc_hd__buf_2 output296 (.A(net296),
    .X(pcpi_rs1[7]));
 sky130_fd_sc_hd__buf_2 output297 (.A(net297),
    .X(pcpi_rs1[8]));
 sky130_fd_sc_hd__buf_2 output298 (.A(net298),
    .X(pcpi_rs1[9]));
 sky130_fd_sc_hd__buf_2 output299 (.A(net299),
    .X(pcpi_rs2[0]));
 sky130_fd_sc_hd__buf_2 output300 (.A(net300),
    .X(pcpi_rs2[10]));
 sky130_fd_sc_hd__buf_2 output301 (.A(net301),
    .X(pcpi_rs2[11]));
 sky130_fd_sc_hd__buf_2 output302 (.A(net302),
    .X(pcpi_rs2[12]));
 sky130_fd_sc_hd__buf_2 output303 (.A(net303),
    .X(pcpi_rs2[13]));
 sky130_fd_sc_hd__buf_2 output304 (.A(net304),
    .X(pcpi_rs2[14]));
 sky130_fd_sc_hd__buf_2 output305 (.A(net305),
    .X(pcpi_rs2[15]));
 sky130_fd_sc_hd__buf_2 output306 (.A(net306),
    .X(pcpi_rs2[16]));
 sky130_fd_sc_hd__buf_2 output307 (.A(net307),
    .X(pcpi_rs2[17]));
 sky130_fd_sc_hd__buf_2 output308 (.A(net308),
    .X(pcpi_rs2[18]));
 sky130_fd_sc_hd__buf_2 output309 (.A(net309),
    .X(pcpi_rs2[19]));
 sky130_fd_sc_hd__buf_2 output310 (.A(net310),
    .X(pcpi_rs2[1]));
 sky130_fd_sc_hd__buf_2 output311 (.A(net311),
    .X(pcpi_rs2[20]));
 sky130_fd_sc_hd__buf_2 output312 (.A(net312),
    .X(pcpi_rs2[21]));
 sky130_fd_sc_hd__buf_2 output313 (.A(net313),
    .X(pcpi_rs2[22]));
 sky130_fd_sc_hd__buf_2 output314 (.A(net314),
    .X(pcpi_rs2[23]));
 sky130_fd_sc_hd__buf_2 output315 (.A(net315),
    .X(pcpi_rs2[24]));
 sky130_fd_sc_hd__buf_2 output316 (.A(net316),
    .X(pcpi_rs2[25]));
 sky130_fd_sc_hd__buf_2 output317 (.A(net317),
    .X(pcpi_rs2[26]));
 sky130_fd_sc_hd__buf_2 output318 (.A(net318),
    .X(pcpi_rs2[27]));
 sky130_fd_sc_hd__buf_2 output319 (.A(net319),
    .X(pcpi_rs2[28]));
 sky130_fd_sc_hd__buf_2 output320 (.A(net320),
    .X(pcpi_rs2[29]));
 sky130_fd_sc_hd__buf_2 output321 (.A(net321),
    .X(pcpi_rs2[2]));
 sky130_fd_sc_hd__buf_2 output322 (.A(net322),
    .X(pcpi_rs2[30]));
 sky130_fd_sc_hd__buf_2 output323 (.A(net323),
    .X(pcpi_rs2[31]));
 sky130_fd_sc_hd__buf_2 output324 (.A(net324),
    .X(pcpi_rs2[3]));
 sky130_fd_sc_hd__buf_2 output325 (.A(net325),
    .X(pcpi_rs2[4]));
 sky130_fd_sc_hd__buf_2 output326 (.A(net326),
    .X(pcpi_rs2[5]));
 sky130_fd_sc_hd__buf_2 output327 (.A(net327),
    .X(pcpi_rs2[6]));
 sky130_fd_sc_hd__buf_2 output328 (.A(net328),
    .X(pcpi_rs2[7]));
 sky130_fd_sc_hd__buf_2 output329 (.A(net329),
    .X(pcpi_rs2[8]));
 sky130_fd_sc_hd__buf_2 output330 (.A(net330),
    .X(pcpi_rs2[9]));
 sky130_fd_sc_hd__clkbuf_4 output331 (.A(net331),
    .X(pcpi_valid));
 sky130_fd_sc_hd__clkbuf_4 output332 (.A(net332),
    .X(trap));
 sky130_fd_sc_hd__buf_1 wire333 (.A(_03347_),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_2 wire334 (.A(_01663_),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_1 max_cap335 (.A(_13793_),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_1 max_cap336 (.A(_12126_),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_1 max_cap337 (.A(_11877_),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_1 max_cap338 (.A(_12001_),
    .X(net338));
 sky130_fd_sc_hd__buf_1 max_cap339 (.A(_12118_),
    .X(net339));
 sky130_fd_sc_hd__buf_1 max_cap340 (.A(_13578_),
    .X(net340));
 sky130_fd_sc_hd__buf_1 max_cap341 (.A(_12653_),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_2 max_cap342 (.A(_12385_),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_1 max_cap343 (.A(_12061_),
    .X(net343));
 sky130_fd_sc_hd__buf_1 wire344 (.A(_13097_),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_1 max_cap345 (.A(net346),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_1 wire346 (.A(_12943_),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_1 max_cap347 (.A(_12651_),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_1 max_cap348 (.A(net349),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_1 wire349 (.A(_13574_),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_1 max_cap350 (.A(_11743_),
    .X(net350));
 sky130_fd_sc_hd__buf_1 max_cap351 (.A(net352),
    .X(net351));
 sky130_fd_sc_hd__buf_1 wire352 (.A(_11524_),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_1 max_cap353 (.A(_11316_),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_1 max_cap354 (.A(_11117_),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_1 max_cap355 (.A(_02048_),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_1 max_cap356 (.A(_01571_),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_1 max_cap357 (.A(net358),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_1 max_cap358 (.A(_11991_),
    .X(net358));
 sky130_fd_sc_hd__buf_1 max_cap359 (.A(_02484_),
    .X(net359));
 sky130_fd_sc_hd__buf_1 max_cap360 (.A(_14065_),
    .X(net360));
 sky130_fd_sc_hd__buf_1 max_cap361 (.A(_13570_),
    .X(net361));
 sky130_fd_sc_hd__buf_1 max_cap362 (.A(_13321_),
    .X(net362));
 sky130_fd_sc_hd__buf_1 max_cap363 (.A(net364),
    .X(net363));
 sky130_fd_sc_hd__buf_1 max_cap364 (.A(_13012_),
    .X(net364));
 sky130_fd_sc_hd__buf_1 max_cap365 (.A(_12729_),
    .X(net365));
 sky130_fd_sc_hd__buf_1 max_cap366 (.A(_13195_),
    .X(net366));
 sky130_fd_sc_hd__buf_1 max_cap367 (.A(_06190_),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_1 wire368 (.A(_08301_),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_2 wire369 (.A(_08225_),
    .X(net369));
 sky130_fd_sc_hd__buf_1 wire370 (.A(_07799_),
    .X(net370));
 sky130_fd_sc_hd__buf_1 wire371 (.A(_10092_),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_2 max_cap372 (.A(_07760_),
    .X(net372));
 sky130_fd_sc_hd__buf_1 max_cap373 (.A(_08223_),
    .X(net373));
 sky130_fd_sc_hd__conb_1 picorv32a_374 (.LO(net374));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_38_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_39_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_40_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_41_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_42_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_43_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_44_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_45_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_46_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_47_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_48_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_49_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_50_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_51_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_52_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_53_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_54_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_55_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_56_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_57_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_58_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_59_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_60_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_61_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_62_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_63_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_64_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_65_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_66_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_67_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_68_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_69_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_70_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_71_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_72_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_73_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_74_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_75_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_76_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_77_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_78_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_79_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_80_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_81_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_82_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_83_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_84_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_85_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_86_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_87_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_88_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_89_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_90_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_91_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_92_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_93_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_94_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_95_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_96_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_97_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_98_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_99_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_100_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_101_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_102_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_103_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_104_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_105_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_106_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_107_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_108_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_109_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_110_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_111_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_112_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_113_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_114_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_115_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_116_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_117_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_118_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_119_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_120_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_121_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_122_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_123_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_124_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_125_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_126_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_127_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_128_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_129_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_130_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_132_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_133_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_134_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_135_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_136_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_137_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_138_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_139_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_140_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_141_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_142_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_143_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_144_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_145_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_146_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_147_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_147_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_148_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_149_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_150_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_151_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_152_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_153_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_153_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_154_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_155_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_156_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_157_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_158_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_158_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_159_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_160_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_160_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_161_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_161_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_162_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_163_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_164_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_165_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_166_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_167_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_168_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_169_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_170_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_171_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_172_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_173_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_174_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_175_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_176_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_177_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_178_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_179_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_180_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_181_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_183_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_184_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_185_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_186_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_187_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_188_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_189_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_189_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_190_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_191_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_192_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_192_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_193_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_193_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_194_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_194_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_195_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_195_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_196_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_197_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_198_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_198_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_200_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_200_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_201_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_201_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_202_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_202_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_203_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_203_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_204_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_204_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_205_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_205_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_207_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_207_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_208_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_208_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_209_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_209_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_210_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_210_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_211_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_211_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_212_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_212_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_213_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_213_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_214_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_214_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_215_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_215_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_216_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_216_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_217_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_217_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_218_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_218_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_219_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_219_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_221_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_221_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_224_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_224_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_225_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_225_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_0__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_1__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_2__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_3__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_4__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_5__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_6__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_7__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_8__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_8__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_9__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_9__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_10__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_10__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_11__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_11__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_12__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_12__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_13__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_13__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_14__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_14__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_15__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_15__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_16__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_16__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_17__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_17__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_18__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_18__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_19__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_19__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_20__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_20__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_21__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_21__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_22__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_22__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_23__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_23__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_24__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_24__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_25__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_25__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_26__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_26__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_27__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_27__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_28__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_28__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_29__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_29__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_30__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_30__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_31__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_31__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload0 (.A(clknet_5_0__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload1 (.A(clknet_5_1__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload2 (.A(clknet_5_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload3 (.A(clknet_5_3__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload4 (.A(clknet_5_4__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload5 (.A(clknet_5_5__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload6 (.A(clknet_5_6__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload7 (.A(clknet_5_9__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload8 (.A(clknet_5_10__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload9 (.A(clknet_5_11__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload10 (.A(clknet_5_12__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload11 (.A(clknet_5_13__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload12 (.A(clknet_5_16__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload13 (.A(clknet_5_17__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload14 (.A(clknet_5_18__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload15 (.A(clknet_5_19__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload16 (.A(clknet_5_20__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload17 (.A(clknet_5_21__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload18 (.A(clknet_5_23__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload19 (.A(clknet_5_24__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload20 (.A(clknet_5_27__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload21 (.A(clknet_5_28__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload22 (.A(clknet_5_29__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload23 (.A(clknet_5_30__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload24 (.A(clknet_5_31__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload25 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__bufinv_16 clkload26 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload27 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__bufinv_16 clkload28 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload29 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload30 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload31 (.A(clknet_leaf_221_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload32 (.A(clknet_leaf_225_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload33 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload34 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload35 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__inv_6 clkload36 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkinv_8 clkload37 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload38 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload39 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload40 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__inv_8 clkload41 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkinv_4 clkload42 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkinv_1 clkload43 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__inv_6 clkload44 (.A(clknet_leaf_213_clk));
 sky130_fd_sc_hd__inv_6 clkload45 (.A(clknet_leaf_217_clk));
 sky130_fd_sc_hd__inv_8 clkload46 (.A(clknet_leaf_219_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload47 (.A(clknet_leaf_214_clk));
 sky130_fd_sc_hd__bufinv_16 clkload48 (.A(clknet_leaf_215_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload49 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload50 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload51 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__bufinv_16 clkload52 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload53 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkinv_4 clkload54 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__inv_6 clkload55 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkinv_4 clkload56 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkinv_4 clkload57 (.A(clknet_leaf_208_clk));
 sky130_fd_sc_hd__inv_6 clkload58 (.A(clknet_leaf_210_clk));
 sky130_fd_sc_hd__inv_6 clkload59 (.A(clknet_leaf_211_clk));
 sky130_fd_sc_hd__inv_6 clkload60 (.A(clknet_leaf_212_clk));
 sky130_fd_sc_hd__inv_8 clkload61 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__bufinv_16 clkload62 (.A(clknet_leaf_42_clk));
 sky130_fd_sc_hd__inv_6 clkload63 (.A(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkinv_4 clkload64 (.A(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload65 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__inv_6 clkload66 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__inv_8 clkload67 (.A(clknet_leaf_53_clk));
 sky130_fd_sc_hd__inv_6 clkload68 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkinv_4 clkload69 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__bufinv_16 clkload70 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkinv_4 clkload71 (.A(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkinv_4 clkload72 (.A(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload73 (.A(clknet_leaf_52_clk));
 sky130_fd_sc_hd__bufinv_16 clkload74 (.A(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload75 (.A(clknet_leaf_55_clk));
 sky130_fd_sc_hd__inv_6 clkload76 (.A(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkinv_4 clkload77 (.A(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload78 (.A(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload79 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__inv_6 clkload80 (.A(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkinv_4 clkload81 (.A(clknet_leaf_59_clk));
 sky130_fd_sc_hd__inv_8 clkload82 (.A(clknet_leaf_60_clk));
 sky130_fd_sc_hd__inv_8 clkload83 (.A(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload84 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkinv_1 clkload85 (.A(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkinv_1 clkload86 (.A(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload87 (.A(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload88 (.A(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkinv_1 clkload89 (.A(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkinv_4 clkload90 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload91 (.A(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkinv_4 clkload92 (.A(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload93 (.A(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkinv_4 clkload94 (.A(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkinv_1 clkload95 (.A(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkinv_4 clkload96 (.A(clknet_leaf_65_clk));
 sky130_fd_sc_hd__bufinv_16 clkload97 (.A(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload98 (.A(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkinv_1 clkload99 (.A(clknet_leaf_71_clk));
 sky130_fd_sc_hd__inv_6 clkload100 (.A(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload101 (.A(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload102 (.A(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkinv_4 clkload103 (.A(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkinv_4 clkload104 (.A(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkinv_1 clkload105 (.A(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload106 (.A(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload107 (.A(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkinv_4 clkload108 (.A(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload109 (.A(clknet_leaf_198_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload110 (.A(clknet_leaf_200_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload111 (.A(clknet_leaf_202_clk));
 sky130_fd_sc_hd__clkinv_4 clkload112 (.A(clknet_leaf_203_clk));
 sky130_fd_sc_hd__inv_6 clkload113 (.A(clknet_leaf_180_clk));
 sky130_fd_sc_hd__inv_6 clkload114 (.A(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkinv_4 clkload115 (.A(clknet_leaf_205_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload116 (.A(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkinv_4 clkload117 (.A(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload118 (.A(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkinv_1 clkload119 (.A(clknet_leaf_207_clk));
 sky130_fd_sc_hd__clkinv_4 clkload120 (.A(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkinv_1 clkload121 (.A(clknet_leaf_172_clk));
 sky130_fd_sc_hd__bufinv_16 clkload122 (.A(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload123 (.A(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload124 (.A(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload125 (.A(clknet_leaf_184_clk));
 sky130_fd_sc_hd__bufinv_16 clkload126 (.A(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload127 (.A(clknet_leaf_186_clk));
 sky130_fd_sc_hd__inv_6 clkload128 (.A(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkinv_4 clkload129 (.A(clknet_leaf_192_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload130 (.A(clknet_leaf_193_clk));
 sky130_fd_sc_hd__clkinv_4 clkload131 (.A(clknet_leaf_194_clk));
 sky130_fd_sc_hd__inv_6 clkload132 (.A(clknet_leaf_195_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload133 (.A(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkinv_4 clkload134 (.A(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload135 (.A(clknet_leaf_158_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload136 (.A(clknet_leaf_159_clk));
 sky130_fd_sc_hd__bufinv_16 clkload137 (.A(clknet_leaf_160_clk));
 sky130_fd_sc_hd__bufinv_16 clkload138 (.A(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkinv_4 clkload139 (.A(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkinv_4 clkload140 (.A(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkinv_4 clkload141 (.A(clknet_leaf_151_clk));
 sky130_fd_sc_hd__inv_6 clkload142 (.A(clknet_leaf_153_clk));
 sky130_fd_sc_hd__bufinv_16 clkload143 (.A(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload144 (.A(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkinv_4 clkload145 (.A(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkinv_1 clkload146 (.A(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkinv_1 clkload147 (.A(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload148 (.A(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload149 (.A(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload150 (.A(clknet_leaf_107_clk));
 sky130_fd_sc_hd__inv_6 clkload151 (.A(clknet_leaf_94_clk));
 sky130_fd_sc_hd__bufinv_16 clkload152 (.A(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload153 (.A(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload154 (.A(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkinv_4 clkload155 (.A(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload156 (.A(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkinv_4 clkload157 (.A(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkinv_4 clkload158 (.A(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload159 (.A(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkinv_4 clkload160 (.A(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload161 (.A(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload162 (.A(clknet_leaf_104_clk));
 sky130_fd_sc_hd__bufinv_16 clkload163 (.A(clknet_leaf_109_clk));
 sky130_fd_sc_hd__inv_6 clkload164 (.A(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload165 (.A(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkinv_4 clkload166 (.A(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkinv_4 clkload167 (.A(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload168 (.A(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkinv_4 clkload169 (.A(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload170 (.A(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkinv_1 clkload171 (.A(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload172 (.A(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkinv_1 clkload173 (.A(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkinv_4 clkload174 (.A(clknet_leaf_119_clk));
 sky130_fd_sc_hd__bufinv_16 clkload175 (.A(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload176 (.A(clknet_leaf_122_clk));
 sky130_fd_sc_hd__bufinv_16 clkload177 (.A(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload178 (.A(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkinv_1 clkload179 (.A(clknet_leaf_161_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload180 (.A(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkinv_4 clkload181 (.A(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload182 (.A(clknet_leaf_143_clk));
 sky130_fd_sc_hd__inv_6 clkload183 (.A(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload184 (.A(clknet_leaf_145_clk));
 sky130_fd_sc_hd__bufinv_16 clkload185 (.A(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkinv_1 clkload186 (.A(clknet_leaf_147_clk));
 sky130_fd_sc_hd__bufinv_16 clkload187 (.A(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload188 (.A(clknet_leaf_149_clk));
 sky130_fd_sc_hd__bufinv_16 clkload189 (.A(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload190 (.A(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkinv_1 clkload191 (.A(clknet_leaf_125_clk));
 sky130_fd_sc_hd__bufinv_16 clkload192 (.A(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkinv_1 clkload193 (.A(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload194 (.A(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload195 (.A(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload196 (.A(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkinv_4 clkload197 (.A(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload198 (.A(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkinv_4 clkload199 (.A(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_1 max_cap1 (.A(_13578_),
    .X(net415));
 sky130_fd_sc_hd__buf_1 max_cap2 (.A(_12653_),
    .X(net416));
 sky130_fd_sc_hd__buf_1 max_cap3 (.A(_13097_),
    .X(net417));
 sky130_fd_sc_hd__buf_1 max_cap4 (.A(_13570_),
    .X(net418));
 sky130_fd_sc_hd__buf_1 max_cap5 (.A(_13012_),
    .X(net419));
 sky130_fd_sc_hd__buf_1 max_cap6 (.A(_12729_),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\alu_add_sub[24] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\alu_add_sub[28] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\alu_out[28] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\alu_add_sub[25] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\alu_add_sub[17] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\alu_add_sub[2] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\alu_add_sub[16] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\alu_add_sub[3] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\alu_add_sub[0] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\alu_add_sub[8] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\alu_add_sub[1] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\alu_add_sub[12] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\alu_add_sub[4] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\alu_add_sub[9] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\alu_add_sub[11] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\alu_add_sub[5] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\alu_add_sub[7] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\alu_add_sub[26] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\alu_add_sub[31] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\irq_mask[9] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\decoded_rd[2] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\alu_add_sub[6] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\alu_add_sub[22] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\decoded_rd[3] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\alu_add_sub[10] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\decoded_rd[1] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(instr_beq),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\irq_mask[10] ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\irq_mask[8] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\alu_add_sub[13] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\decoded_rd[0] ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\irq_mask[12] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(instr_addi),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\mem_rdata_q[28] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\alu_add_sub[14] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(instr_srli),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(instr_add),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\irq_mask[11] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\mem_wordsize[0] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\alu_add_sub[19] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\alu_add_sub[20] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\alu_add_sub[27] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\alu_add_sub[29] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(instr_xori),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\alu_add_sub[15] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\pcpi_timeout_counter[3] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(instr_srl),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(instr_bltu),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(instr_rdcycle),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(instr_and),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(instr_andi),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(instr_slti),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(instr_sltu),
    .X(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_00037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_00037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_00078_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_00078_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_00078_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_00078_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_00078_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_00079_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_00079_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_00079_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_00079_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_00079_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_00079_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_00079_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_00079_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_00079_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_00081_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_00081_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_00081_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_00081_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_00081_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_00082_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_00082_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_00084_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_00084_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_00088_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_00088_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_00088_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_00088_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_00089_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_00090_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_00090_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_00093_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_00096_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_00100_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_00621_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_00725_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_01066_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_01547_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_01547_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_01547_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_01547_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_01547_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_01583_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_01625_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_02147_));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_02147_));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_03633_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_04254_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_04254_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_04755_));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(_05068_));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(_05094_));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(_05145_));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(_05181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(_05181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(_05181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(_05181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(_05182_));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(_05205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(_05205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(_05205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(_05205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(_05302_));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(_05302_));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(_05308_));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(_05542_));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(_05544_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(_05546_));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(_05686_));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(_05686_));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(_05694_));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(_05714_));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(_05714_));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(_05718_));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(_06180_));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(_06302_));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(_07035_));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(_07105_));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(_07388_));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(_07693_));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(_08176_));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(_08176_));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(_08224_));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(_08309_));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(_08309_));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(_08322_));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(_08332_));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(_08338_));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(_08359_));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(_08412_));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(_08412_));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(_08412_));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(_08427_));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(_08436_));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(_08505_));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(_08520_));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(_08525_));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(_08536_));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(_08593_));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(_08696_));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(_08736_));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(_08798_));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(_08978_));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(_09091_));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(_09149_));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(_09319_));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(_09339_));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(_09420_));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(_09590_));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(_09626_));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(_09626_));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(_09626_));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(_09704_));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(_09704_));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(_09704_));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(_09739_));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(_09744_));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(_09744_));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(_09781_));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(_09855_));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(_09966_));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(_10003_));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(_10197_));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(_10197_));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(_10197_));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(_10206_));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(_10206_));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(_10214_));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(_10224_));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(_10241_));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(_10246_));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(_10250_));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(_10250_));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(_10264_));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(_10264_));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(_10273_));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(_10277_));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(_10279_));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(_10331_));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(_10334_));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(_10334_));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(_10354_));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(_10354_));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(_10367_));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(_10372_));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(_10378_));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(_10378_));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(_10389_));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(_10389_));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(_10389_));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(_10392_));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(_10392_));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(_10600_));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(_10603_));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(_10609_));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(_10738_));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(_10760_));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(_10760_));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(_10784_));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(_10788_));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(_10958_));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(_10964_));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(_11048_));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(_11109_));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(_11137_));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(_11137_));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(_11137_));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(_11142_));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(_11157_));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(_11157_));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(_11157_));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(_11167_));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(_11201_));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(_11201_));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(_11201_));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(_11237_));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(_11237_));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(_11237_));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(_11237_));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(_11264_));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(_11265_));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(_11277_));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(_11297_));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(_11353_));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(_11353_));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(_11353_));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(_11353_));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(_11368_));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(_11447_));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(_11447_));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(_11474_));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(_11482_));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(_11482_));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(_11590_));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(_11590_));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(_11662_));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(_11662_));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(_11666_));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(_11707_));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(_11773_));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(_11826_));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(_11831_));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(_11958_));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(_11961_));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(_11961_));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(_12044_));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(_12044_));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(_12067_));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(_12067_));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(_12098_));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(_12146_));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(_12282_));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(_12282_));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(_12282_));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(_12282_));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(_12325_));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(_12586_));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(_12586_));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(_13057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(_13228_));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(_13228_));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(_13442_));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(_13442_));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(_13447_));
 sky130_fd_sc_hd__diode_2 ANTENNA_268 (.DIODE(_13447_));
 sky130_fd_sc_hd__diode_2 ANTENNA_269 (.DIODE(_13754_));
 sky130_fd_sc_hd__diode_2 ANTENNA_270 (.DIODE(_13819_));
 sky130_fd_sc_hd__diode_2 ANTENNA_271 (.DIODE(_13820_));
 sky130_fd_sc_hd__diode_2 ANTENNA_272 (.DIODE(_13820_));
 sky130_fd_sc_hd__diode_2 ANTENNA_273 (.DIODE(_13821_));
 sky130_fd_sc_hd__diode_2 ANTENNA_274 (.DIODE(_13821_));
 sky130_fd_sc_hd__diode_2 ANTENNA_275 (.DIODE(_13849_));
 sky130_fd_sc_hd__diode_2 ANTENNA_276 (.DIODE(_13849_));
 sky130_fd_sc_hd__diode_2 ANTENNA_277 (.DIODE(_13858_));
 sky130_fd_sc_hd__diode_2 ANTENNA_278 (.DIODE(_13858_));
 sky130_fd_sc_hd__diode_2 ANTENNA_279 (.DIODE(_13901_));
 sky130_fd_sc_hd__diode_2 ANTENNA_280 (.DIODE(_14105_));
 sky130_fd_sc_hd__diode_2 ANTENNA_281 (.DIODE(_14283_));
 sky130_fd_sc_hd__diode_2 ANTENNA_282 (.DIODE(\alu_out[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_283 (.DIODE(\alu_out[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_284 (.DIODE(\alu_out_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_285 (.DIODE(\alu_out_q[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_286 (.DIODE(\alu_out_q[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_287 (.DIODE(\alu_out_q[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_288 (.DIODE(\alu_out_q[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_289 (.DIODE(\alu_out_q[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_290 (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_291 (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_292 (.DIODE(\decoded_imm[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_293 (.DIODE(\decoded_imm_uj[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_294 (.DIODE(\decoded_imm_uj[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_295 (.DIODE(\genblk1.pcpi_mul.rd[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_296 (.DIODE(\genblk1.pcpi_mul.rd[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_297 (.DIODE(\genblk1.pcpi_mul.rd[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_298 (.DIODE(\genblk1.pcpi_mul.rd[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_299 (.DIODE(\genblk1.pcpi_mul.rd[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_300 (.DIODE(\genblk1.pcpi_mul.rd[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_301 (.DIODE(\genblk1.pcpi_mul.rd[50] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_302 (.DIODE(\genblk1.pcpi_mul.rd[58] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_303 (.DIODE(\genblk1.pcpi_mul.rd[58] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_304 (.DIODE(\genblk1.pcpi_mul.rd[58] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_305 (.DIODE(\genblk1.pcpi_mul.rd[58] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_306 (.DIODE(\genblk1.pcpi_mul.rd[58] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_307 (.DIODE(\genblk1.pcpi_mul.rd[58] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_308 (.DIODE(\genblk1.pcpi_mul.rd[58] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_309 (.DIODE(\genblk1.pcpi_mul.rd[58] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_310 (.DIODE(\genblk1.pcpi_mul.rd[59] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_311 (.DIODE(\genblk1.pcpi_mul.rd[59] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_312 (.DIODE(\genblk1.pcpi_mul.rd[59] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_313 (.DIODE(\genblk1.pcpi_mul.rd[59] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_314 (.DIODE(\genblk1.pcpi_mul.rd[59] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_315 (.DIODE(\genblk1.pcpi_mul.rd[59] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_316 (.DIODE(\genblk1.pcpi_mul.rd[59] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_317 (.DIODE(\genblk1.pcpi_mul.rd[59] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_318 (.DIODE(\genblk1.pcpi_mul.rd[59] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_319 (.DIODE(\genblk1.pcpi_mul.rd[59] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_320 (.DIODE(\genblk1.pcpi_mul.rd[61] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_321 (.DIODE(\genblk1.pcpi_mul.rd[61] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_322 (.DIODE(\genblk1.pcpi_mul.rd[61] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_323 (.DIODE(\genblk1.pcpi_mul.rd[61] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_324 (.DIODE(\genblk1.pcpi_mul.rd[61] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_325 (.DIODE(\genblk1.pcpi_mul.rd[61] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_326 (.DIODE(\genblk1.pcpi_mul.rd[61] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_327 (.DIODE(\genblk1.pcpi_mul.rd[61] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_328 (.DIODE(\genblk1.pcpi_mul.rd[62] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_329 (.DIODE(\genblk1.pcpi_mul.rd[62] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_330 (.DIODE(\genblk1.pcpi_mul.rd[62] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_331 (.DIODE(\genblk1.pcpi_mul.rd[62] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_332 (.DIODE(\genblk1.pcpi_mul.rd[62] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_333 (.DIODE(\genblk1.pcpi_mul.rd[62] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_334 (.DIODE(\genblk1.pcpi_mul.rd[62] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_335 (.DIODE(\genblk1.pcpi_mul.rd[62] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_336 (.DIODE(\genblk1.pcpi_mul.rd[63] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_337 (.DIODE(\genblk1.pcpi_mul.rd[63] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_338 (.DIODE(\genblk1.pcpi_mul.rd[63] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_339 (.DIODE(\genblk1.pcpi_mul.rd[63] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_340 (.DIODE(\genblk1.pcpi_mul.rd[63] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_341 (.DIODE(\genblk1.pcpi_mul.rd[63] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_342 (.DIODE(\genblk1.pcpi_mul.rs1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_343 (.DIODE(\genblk1.pcpi_mul.rs1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_344 (.DIODE(\genblk1.pcpi_mul.rs1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_345 (.DIODE(\genblk1.pcpi_mul.rs1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_346 (.DIODE(\genblk1.pcpi_mul.rs1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_347 (.DIODE(\genblk1.pcpi_mul.rs1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_348 (.DIODE(\genblk1.pcpi_mul.rs2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_349 (.DIODE(\genblk1.pcpi_mul.rs2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_350 (.DIODE(\mem_rdata_q[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_351 (.DIODE(\mem_rdata_q[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_352 (.DIODE(\mem_rdata_q[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_353 (.DIODE(\reg_next_pc[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_354 (.DIODE(\reg_next_pc[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_355 (.DIODE(\reg_next_pc[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_356 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_357 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_358 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_359 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_360 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_361 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_362 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_363 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_364 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_365 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_366 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_367 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_368 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_369 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_370 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_371 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_372 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_373 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_374 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_375 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_376 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_377 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_378 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_379 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_380 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_381 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_382 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_383 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_384 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_385 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_386 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_387 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_388 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_389 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_390 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_391 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_392 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_393 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_394 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_395 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_396 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_397 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_398 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_399 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_400 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_401 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_402 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_403 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_404 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_405 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_406 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_407 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_408 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_409 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_410 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_411 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_412 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_413 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_414 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_415 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_416 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_417 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_418 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_419 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_420 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_421 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_422 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_423 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_424 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_425 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_426 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_427 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_428 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_429 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_430 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_431 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_432 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_433 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_434 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_435 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_436 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_437 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_438 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_439 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_440 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_441 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_442 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_443 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_444 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_445 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_446 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_447 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_448 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_449 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_450 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_451 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_452 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_453 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_454 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_455 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_456 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_457 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_458 (.DIODE(_00097_));
 sky130_fd_sc_hd__diode_2 ANTENNA_459 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA_460 (.DIODE(_02713_));
 sky130_fd_sc_hd__diode_2 ANTENNA_461 (.DIODE(_04988_));
 sky130_fd_sc_hd__diode_2 ANTENNA_462 (.DIODE(_05172_));
 sky130_fd_sc_hd__diode_2 ANTENNA_463 (.DIODE(_05172_));
 sky130_fd_sc_hd__diode_2 ANTENNA_464 (.DIODE(_08412_));
 sky130_fd_sc_hd__diode_2 ANTENNA_465 (.DIODE(_08412_));
 sky130_fd_sc_hd__diode_2 ANTENNA_466 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_467 (.DIODE(_09205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_468 (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA_469 (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA_470 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_471 (.DIODE(_09590_));
 sky130_fd_sc_hd__diode_2 ANTENNA_472 (.DIODE(_09626_));
 sky130_fd_sc_hd__diode_2 ANTENNA_473 (.DIODE(_09667_));
 sky130_fd_sc_hd__diode_2 ANTENNA_474 (.DIODE(_09667_));
 sky130_fd_sc_hd__diode_2 ANTENNA_475 (.DIODE(_10108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_476 (.DIODE(_10108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_477 (.DIODE(_10108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_478 (.DIODE(_10108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_479 (.DIODE(_10108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_480 (.DIODE(_10108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_481 (.DIODE(_10108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_482 (.DIODE(_10108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_483 (.DIODE(_10108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_484 (.DIODE(_10108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_485 (.DIODE(_10108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_486 (.DIODE(_10108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_487 (.DIODE(_10108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_488 (.DIODE(_10108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_489 (.DIODE(_10108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_490 (.DIODE(_10108_));
 sky130_fd_sc_hd__diode_2 ANTENNA_491 (.DIODE(_10157_));
 sky130_fd_sc_hd__diode_2 ANTENNA_492 (.DIODE(_10157_));
 sky130_fd_sc_hd__diode_2 ANTENNA_493 (.DIODE(_10157_));
 sky130_fd_sc_hd__diode_2 ANTENNA_494 (.DIODE(_10255_));
 sky130_fd_sc_hd__diode_2 ANTENNA_495 (.DIODE(_10736_));
 sky130_fd_sc_hd__diode_2 ANTENNA_496 (.DIODE(_11369_));
 sky130_fd_sc_hd__diode_2 ANTENNA_497 (.DIODE(_11481_));
 sky130_fd_sc_hd__diode_2 ANTENNA_498 (.DIODE(_11949_));
 sky130_fd_sc_hd__diode_2 ANTENNA_499 (.DIODE(_11949_));
 sky130_fd_sc_hd__diode_2 ANTENNA_500 (.DIODE(_11949_));
 sky130_fd_sc_hd__diode_2 ANTENNA_501 (.DIODE(_11961_));
 sky130_fd_sc_hd__diode_2 ANTENNA_502 (.DIODE(_13614_));
 sky130_fd_sc_hd__diode_2 ANTENNA_503 (.DIODE(_13614_));
 sky130_fd_sc_hd__diode_2 ANTENNA_504 (.DIODE(\genblk1.pcpi_mul.rd[60] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_505 (.DIODE(\genblk1.pcpi_mul.rs1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_506 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_507 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_508 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_509 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_510 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_511 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_512 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_513 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_514 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_515 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_516 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_517 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_518 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_519 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_520 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_521 (.DIODE(_00089_));
 sky130_fd_sc_hd__diode_2 ANTENNA_522 (.DIODE(_00089_));
 sky130_fd_sc_hd__diode_2 ANTENNA_523 (.DIODE(_00089_));
 sky130_fd_sc_hd__diode_2 ANTENNA_524 (.DIODE(_09245_));
 sky130_fd_sc_hd__diode_2 ANTENNA_525 (.DIODE(_09245_));
 sky130_fd_sc_hd__diode_2 ANTENNA_526 (.DIODE(_10003_));
 sky130_fd_sc_hd__diode_2 ANTENNA_527 (.DIODE(\genblk1.pcpi_mul.rd[49] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_528 (.DIODE(_00089_));
 sky130_fd_sc_hd__diode_2 ANTENNA_529 (.DIODE(_00089_));
 sky130_fd_sc_hd__diode_2 ANTENNA_530 (.DIODE(_00089_));
 sky130_fd_sc_hd__diode_2 ANTENNA_531 (.DIODE(_00089_));
 sky130_fd_sc_hd__diode_2 ANTENNA_532 (.DIODE(_00089_));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1064 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_926 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1094 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_983 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_924 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_947 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1066 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1226 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1098 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_870 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1392 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1092 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1008 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_927 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_898 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1059 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1098 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1038 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1066 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1074 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1043 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1422 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_1472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1450 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_1410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1092 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1094 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_926 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1043 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1092 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_1453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_1312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_1409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_1298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_1409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_1376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_868 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1043 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1066 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_1324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_1421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_1410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_1397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_1446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_1382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_1424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_1429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_1468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1036 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_1327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_1292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_871 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_1310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_1366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_1429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_1442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_1371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_1389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_927 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_1290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_1370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_1394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_1468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_1392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213_1407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_1435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_213_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_1250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_214_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_1358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_1384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_1397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_1179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216_1402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_1474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_1310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_1380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_219_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_1208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_1372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_219_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_1408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_952 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_222_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_222_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_222_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_222_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_222_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_222_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_222_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_222_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_222_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_222_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_954 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_222_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_222_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_222_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_223_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_223_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_223_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_223_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_223_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_223_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_223_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_1448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_224_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_224_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_224_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_224_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_224_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_224_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_224_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_224_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_224_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_224_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_896 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_224_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_224_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_224_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_224_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_224_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_224_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_224_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_224_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_1389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_224_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_224_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_1336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_1199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_230_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_230_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_230_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_230_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_230_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_230_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_230_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_230_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_230_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_230_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_230_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_230_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_230_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_1314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230_1326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_230_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_230_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_231_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_231_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_231_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_231_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_231_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_231_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_231_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_231_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_231_1208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_231_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_231_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_232_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_232_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_232_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_232_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_232_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_232_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_232_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_232_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_232_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_232_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_232_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_232_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_232_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_232_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_232_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_232_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_232_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_232_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_232_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_232_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_232_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_232_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_232_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_232_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_232_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_232_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_232_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_232_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_232_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_232_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_232_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_232_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_232_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_232_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_233_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_233_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_233_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_233_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_233_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_234_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_234_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_234_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_234_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_234_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_234_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_234_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_234_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_234_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_234_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_234_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_234_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_234_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_234_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_234_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_234_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_234_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_234_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_234_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_234_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_234_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_234_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_234_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_234_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_234_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_234_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_234_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_234_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_235_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_235_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_235_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_235_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_235_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_235_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_235_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_235_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_235_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_235_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_235_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_235_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_235_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_235_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_235_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_235_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_235_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_235_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_235_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_235_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_235_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_235_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_235_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_235_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1098 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_235_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_235_1148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_235_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_235_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_235_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_235_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_235_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_235_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_236_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_236_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_236_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_236_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_236_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_236_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_236_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_236_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_236_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_236_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_236_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_236_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_236_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_236_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_236_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_236_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_236_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_236_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_236_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_236_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_236_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_236_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_236_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_236_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_236_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_236_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_236_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_236_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_236_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_236_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_236_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_237_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_237_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_237_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_237_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_237_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_237_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_237_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_237_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_237_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_237_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_237_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_237_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_237_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_237_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_237_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_237_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_237_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_237_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_237_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_237_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_237_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_237_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_1264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_237_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_1277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_237_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_237_1316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_237_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_238_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_238_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_238_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_238_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_238_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_238_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_238_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_238_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_238_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_238_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_238_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_238_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_238_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_238_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_238_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_238_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_238_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_238_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_238_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_238_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_238_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_238_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_238_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_238_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_238_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_238_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_238_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_238_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_238_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_238_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_238_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_238_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_238_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_238_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_238_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_239_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_239_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_239_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_239_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_239_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_239_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_239_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_239_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_239_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_239_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_239_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_239_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_239_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_1299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_239_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_240_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_240_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_240_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_240_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_240_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_240_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_240_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_240_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_240_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_240_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_240_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_240_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_240_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_240_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_240_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_240_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_240_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_240_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_240_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_240_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_240_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_240_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_240_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_240_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_240_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_240_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_240_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_240_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_240_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_240_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_240_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_240_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_240_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_240_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_240_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_240_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_240_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_240_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_240_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_240_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_240_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_240_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_240_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_240_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_240_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_240_1278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_240_1303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_240_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_240_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_240_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_241_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_241_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_241_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_241_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_241_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_241_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_241_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_241_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_241_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_241_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_241_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_241_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_241_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_241_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_241_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_241_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_241_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_241_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_241_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_241_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_241_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_241_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_241_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_241_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_241_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_241_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_241_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_241_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_241_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_241_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_241_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_241_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_241_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_241_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_241_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_241_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_241_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_242_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_242_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_242_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_242_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_242_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_242_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_242_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_242_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_242_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_242_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_242_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_242_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_242_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_242_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_242_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_242_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_242_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_242_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_242_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_242_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_242_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_242_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_242_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_242_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_242_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_242_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_242_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_242_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_242_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_242_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_242_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_242_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_242_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_243_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_243_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_243_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_243_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_243_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_243_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_243_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_243_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_243_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_243_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_243_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_243_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243_1152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_243_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_244_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_244_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_244_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_244_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_244_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_244_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_244_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_244_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_244_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_244_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_244_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_244_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_244_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_244_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_244_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_244_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_244_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_244_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_244_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_244_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_244_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_244_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_244_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_244_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_245_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_245_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_245_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_245_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_245_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_245_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_245_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_245_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_245_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_245_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_245_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_245_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_245_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_245_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_245_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_245_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_245_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_245_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_246_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_246_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_246_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_246_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_246_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_246_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_246_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_246_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_246_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_246_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_246_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_246_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_246_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_246_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_246_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_246_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_246_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_246_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_246_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_246_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_246_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_246_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_246_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_246_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_246_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_246_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_246_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_246_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_246_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_246_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_246_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_247_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_247_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_247_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_247_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_247_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_247_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_247_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_247_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_247_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_247_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_247_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_247_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_247_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_247_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_247_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_247_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_247_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_247_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_247_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_247_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_247_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_247_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_247_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_247_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_247_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_247_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_248_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_248_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_248_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_248_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_248_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_248_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_248_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_248_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_248_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_248_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_248_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_248_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_248_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_248_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_248_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_248_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_248_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_248_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_248_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_248_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_248_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_248_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_248_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_248_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_248_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_248_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_248_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_248_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_248_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_248_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_248_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_248_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_248_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_248_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_248_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_248_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_248_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_248_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_248_1473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_249_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1043 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1469 ();
 assign mem_addr[0] = net374;
 assign mem_addr[1] = net375;
 assign mem_la_addr[0] = net376;
 assign mem_la_addr[1] = net377;
 assign trace_data[0] = net378;
 assign trace_data[10] = net388;
 assign trace_data[11] = net389;
 assign trace_data[12] = net390;
 assign trace_data[13] = net391;
 assign trace_data[14] = net392;
 assign trace_data[15] = net393;
 assign trace_data[16] = net394;
 assign trace_data[17] = net395;
 assign trace_data[18] = net396;
 assign trace_data[19] = net397;
 assign trace_data[1] = net379;
 assign trace_data[20] = net398;
 assign trace_data[21] = net399;
 assign trace_data[22] = net400;
 assign trace_data[23] = net401;
 assign trace_data[24] = net402;
 assign trace_data[25] = net403;
 assign trace_data[26] = net404;
 assign trace_data[27] = net405;
 assign trace_data[28] = net406;
 assign trace_data[29] = net407;
 assign trace_data[2] = net380;
 assign trace_data[30] = net408;
 assign trace_data[31] = net409;
 assign trace_data[32] = net410;
 assign trace_data[33] = net411;
 assign trace_data[34] = net412;
 assign trace_data[35] = net413;
 assign trace_data[3] = net381;
 assign trace_data[4] = net382;
 assign trace_data[5] = net383;
 assign trace_data[6] = net384;
 assign trace_data[7] = net385;
 assign trace_data[8] = net386;
 assign trace_data[9] = net387;
 assign trace_valid = net414;
endmodule
